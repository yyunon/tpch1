-------------------------------------
-- Defines the dataPath width
--
-------------------------------------
package mypackage is
   constant XBITS :INTEGER := 64; 
   constant YBITS :INTEGER := 64;
   constant GRAIN :INTEGER := 2; --Allways in 2!!!!
   constant DEPTH :INTEGER := 4; --Every how much steps register
end mypackage;
