-- Copyright 2018-2019 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
-- This file was generated by Fletchgen. Modify this file at your own risk.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.Array_pkg.all;

entity PriceSummaryWriter_l is
  generic (
    INDEX_WIDTH                         : integer := 32;
    TAG_WIDTH                           : integer := 1;
    L_RETURNFLAG_O_BUS_ADDR_WIDTH       : integer := 64;
    L_RETURNFLAG_O_BUS_DATA_WIDTH       : integer := 512;
    L_RETURNFLAG_O_BUS_LEN_WIDTH        : integer := 8;
    L_RETURNFLAG_O_BUS_BURST_STEP_LEN   : integer := 1;
    L_RETURNFLAG_O_BUS_BURST_MAX_LEN    : integer := 16;
    L_LINESTATUS_O_BUS_ADDR_WIDTH       : integer := 64;
    L_LINESTATUS_O_BUS_DATA_WIDTH       : integer := 512;
    L_LINESTATUS_O_BUS_LEN_WIDTH        : integer := 8;
    L_LINESTATUS_O_BUS_BURST_STEP_LEN   : integer := 1;
    L_LINESTATUS_O_BUS_BURST_MAX_LEN    : integer := 16;
    L_SUM_QTY_BUS_ADDR_WIDTH            : integer := 64;
    L_SUM_QTY_BUS_DATA_WIDTH            : integer := 512;
    L_SUM_QTY_BUS_LEN_WIDTH             : integer := 8;
    L_SUM_QTY_BUS_BURST_STEP_LEN        : integer := 1;
    L_SUM_QTY_BUS_BURST_MAX_LEN         : integer := 16;
    L_SUM_BASE_PRICE_BUS_ADDR_WIDTH     : integer := 64;
    L_SUM_BASE_PRICE_BUS_DATA_WIDTH     : integer := 512;
    L_SUM_BASE_PRICE_BUS_LEN_WIDTH      : integer := 8;
    L_SUM_BASE_PRICE_BUS_BURST_STEP_LEN : integer := 1;
    L_SUM_BASE_PRICE_BUS_BURST_MAX_LEN  : integer := 16;
    L_SUM_DISC_PRICE_BUS_ADDR_WIDTH     : integer := 64;
    L_SUM_DISC_PRICE_BUS_DATA_WIDTH     : integer := 512;
    L_SUM_DISC_PRICE_BUS_LEN_WIDTH      : integer := 8;
    L_SUM_DISC_PRICE_BUS_BURST_STEP_LEN : integer := 1;
    L_SUM_DISC_PRICE_BUS_BURST_MAX_LEN  : integer := 16;
    L_SUM_CHARGE_BUS_ADDR_WIDTH         : integer := 64;
    L_SUM_CHARGE_BUS_DATA_WIDTH         : integer := 512;
    L_SUM_CHARGE_BUS_LEN_WIDTH          : integer := 8;
    L_SUM_CHARGE_BUS_BURST_STEP_LEN     : integer := 1;
    L_SUM_CHARGE_BUS_BURST_MAX_LEN      : integer := 16;
    L_AVG_QTY_BUS_ADDR_WIDTH            : integer := 64;
    L_AVG_QTY_BUS_DATA_WIDTH            : integer := 512;
    L_AVG_QTY_BUS_LEN_WIDTH             : integer := 8;
    L_AVG_QTY_BUS_BURST_STEP_LEN        : integer := 1;
    L_AVG_QTY_BUS_BURST_MAX_LEN         : integer := 16;
    L_AVG_PRICE_BUS_ADDR_WIDTH          : integer := 64;
    L_AVG_PRICE_BUS_DATA_WIDTH          : integer := 512;
    L_AVG_PRICE_BUS_LEN_WIDTH           : integer := 8;
    L_AVG_PRICE_BUS_BURST_STEP_LEN      : integer := 1;
    L_AVG_PRICE_BUS_BURST_MAX_LEN       : integer := 16;
    L_AVG_DISC_BUS_ADDR_WIDTH           : integer := 64;
    L_AVG_DISC_BUS_DATA_WIDTH           : integer := 512;
    L_AVG_DISC_BUS_LEN_WIDTH            : integer := 8;
    L_AVG_DISC_BUS_BURST_STEP_LEN       : integer := 1;
    L_AVG_DISC_BUS_BURST_MAX_LEN        : integer := 16;
    L_COUNT_ORDER_BUS_ADDR_WIDTH        : integer := 64;
    L_COUNT_ORDER_BUS_DATA_WIDTH        : integer := 512;
    L_COUNT_ORDER_BUS_LEN_WIDTH         : integer := 8;
    L_COUNT_ORDER_BUS_BURST_STEP_LEN    : integer := 1;
    L_COUNT_ORDER_BUS_BURST_MAX_LEN     : integer := 16
  );
  port (
    bcd_clk                          : in  std_logic;
    bcd_reset                        : in  std_logic;
    kcd_clk                          : in  std_logic;
    kcd_reset                        : in  std_logic;
    l_returnflag_o_valid             : in  std_logic;
    l_returnflag_o_ready             : out std_logic;
    l_returnflag_o_dvalid            : in  std_logic;
    l_returnflag_o_last              : in  std_logic;
    l_returnflag_o_length            : in  std_logic_vector(31 downto 0);
    l_returnflag_o_count             : in  std_logic_vector(0 downto 0);
    l_returnflag_o_chars_valid       : in  std_logic;
    l_returnflag_o_chars_ready       : out std_logic;
    l_returnflag_o_chars_dvalid      : in  std_logic;
    l_returnflag_o_chars_last        : in  std_logic;
    l_returnflag_o_chars             : in  std_logic_vector(7 downto 0);
    l_returnflag_o_chars_count       : in  std_logic_vector(0 downto 0);
    l_returnflag_o_bus_wreq_valid    : out std_logic;
    l_returnflag_o_bus_wreq_ready    : in  std_logic;
    l_returnflag_o_bus_wreq_addr     : out std_logic_vector(L_RETURNFLAG_O_BUS_ADDR_WIDTH-1 downto 0);
    l_returnflag_o_bus_wreq_len      : out std_logic_vector(L_RETURNFLAG_O_BUS_LEN_WIDTH-1 downto 0);
    l_returnflag_o_bus_wdat_valid    : out std_logic;
    l_returnflag_o_bus_wdat_ready    : in  std_logic;
    l_returnflag_o_bus_wdat_data     : out std_logic_vector(L_RETURNFLAG_O_BUS_DATA_WIDTH-1 downto 0);
    l_returnflag_o_bus_wdat_strobe   : out std_logic_vector(L_RETURNFLAG_O_BUS_DATA_WIDTH/8-1 downto 0);
    l_returnflag_o_bus_wdat_last     : out std_logic;
    l_returnflag_o_cmd_valid         : in  std_logic;
    l_returnflag_o_cmd_ready         : out std_logic;
    l_returnflag_o_cmd_firstIdx      : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_returnflag_o_cmd_lastIdx       : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_returnflag_o_cmd_ctrl          : in  std_logic_vector(L_RETURNFLAG_O_BUS_ADDR_WIDTH*2-1 downto 0);
    l_returnflag_o_cmd_tag           : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_returnflag_o_unl_valid         : out std_logic;
    l_returnflag_o_unl_ready         : in  std_logic;
    l_returnflag_o_unl_tag           : out std_logic_vector(TAG_WIDTH-1 downto 0);
    l_linestatus_o_valid             : in  std_logic;
    l_linestatus_o_ready             : out std_logic;
    l_linestatus_o_dvalid            : in  std_logic;
    l_linestatus_o_last              : in  std_logic;
    l_linestatus_o_length            : in  std_logic_vector(31 downto 0);
    l_linestatus_o_count             : in  std_logic_vector(0 downto 0);
    l_linestatus_o_chars_valid       : in  std_logic;
    l_linestatus_o_chars_ready       : out std_logic;
    l_linestatus_o_chars_dvalid      : in  std_logic;
    l_linestatus_o_chars_last        : in  std_logic;
    l_linestatus_o_chars             : in  std_logic_vector(7 downto 0);
    l_linestatus_o_chars_count       : in  std_logic_vector(0 downto 0);
    l_linestatus_o_bus_wreq_valid    : out std_logic;
    l_linestatus_o_bus_wreq_ready    : in  std_logic;
    l_linestatus_o_bus_wreq_addr     : out std_logic_vector(L_LINESTATUS_O_BUS_ADDR_WIDTH-1 downto 0);
    l_linestatus_o_bus_wreq_len      : out std_logic_vector(L_LINESTATUS_O_BUS_LEN_WIDTH-1 downto 0);
    l_linestatus_o_bus_wdat_valid    : out std_logic;
    l_linestatus_o_bus_wdat_ready    : in  std_logic;
    l_linestatus_o_bus_wdat_data     : out std_logic_vector(L_LINESTATUS_O_BUS_DATA_WIDTH-1 downto 0);
    l_linestatus_o_bus_wdat_strobe   : out std_logic_vector(L_LINESTATUS_O_BUS_DATA_WIDTH/8-1 downto 0);
    l_linestatus_o_bus_wdat_last     : out std_logic;
    l_linestatus_o_cmd_valid         : in  std_logic;
    l_linestatus_o_cmd_ready         : out std_logic;
    l_linestatus_o_cmd_firstIdx      : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_linestatus_o_cmd_lastIdx       : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_linestatus_o_cmd_ctrl          : in  std_logic_vector(L_LINESTATUS_O_BUS_ADDR_WIDTH*2-1 downto 0);
    l_linestatus_o_cmd_tag           : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_linestatus_o_unl_valid         : out std_logic;
    l_linestatus_o_unl_ready         : in  std_logic;
    l_linestatus_o_unl_tag           : out std_logic_vector(TAG_WIDTH-1 downto 0);
    l_sum_qty_valid                  : in  std_logic;
    l_sum_qty_ready                  : out std_logic;
    l_sum_qty_dvalid                 : in  std_logic;
    l_sum_qty_last                   : in  std_logic;
    l_sum_qty                        : in  std_logic_vector(63 downto 0);
    l_sum_qty_bus_wreq_valid         : out std_logic;
    l_sum_qty_bus_wreq_ready         : in  std_logic;
    l_sum_qty_bus_wreq_addr          : out std_logic_vector(L_SUM_QTY_BUS_ADDR_WIDTH-1 downto 0);
    l_sum_qty_bus_wreq_len           : out std_logic_vector(L_SUM_QTY_BUS_LEN_WIDTH-1 downto 0);
    l_sum_qty_bus_wdat_valid         : out std_logic;
    l_sum_qty_bus_wdat_ready         : in  std_logic;
    l_sum_qty_bus_wdat_data          : out std_logic_vector(L_SUM_QTY_BUS_DATA_WIDTH-1 downto 0);
    l_sum_qty_bus_wdat_strobe        : out std_logic_vector(L_SUM_QTY_BUS_DATA_WIDTH/8-1 downto 0);
    l_sum_qty_bus_wdat_last          : out std_logic;
    l_sum_qty_cmd_valid              : in  std_logic;
    l_sum_qty_cmd_ready              : out std_logic;
    l_sum_qty_cmd_firstIdx           : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_sum_qty_cmd_lastIdx            : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_sum_qty_cmd_ctrl               : in  std_logic_vector(L_SUM_QTY_BUS_ADDR_WIDTH-1 downto 0);
    l_sum_qty_cmd_tag                : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_sum_qty_unl_valid              : out std_logic;
    l_sum_qty_unl_ready              : in  std_logic;
    l_sum_qty_unl_tag                : out std_logic_vector(TAG_WIDTH-1 downto 0);
    l_sum_base_price_valid           : in  std_logic;
    l_sum_base_price_ready           : out std_logic;
    l_sum_base_price_dvalid          : in  std_logic;
    l_sum_base_price_last            : in  std_logic;
    l_sum_base_price                 : in  std_logic_vector(63 downto 0);
    l_sum_base_price_bus_wreq_valid  : out std_logic;
    l_sum_base_price_bus_wreq_ready  : in  std_logic;
    l_sum_base_price_bus_wreq_addr   : out std_logic_vector(L_SUM_BASE_PRICE_BUS_ADDR_WIDTH-1 downto 0);
    l_sum_base_price_bus_wreq_len    : out std_logic_vector(L_SUM_BASE_PRICE_BUS_LEN_WIDTH-1 downto 0);
    l_sum_base_price_bus_wdat_valid  : out std_logic;
    l_sum_base_price_bus_wdat_ready  : in  std_logic;
    l_sum_base_price_bus_wdat_data   : out std_logic_vector(L_SUM_BASE_PRICE_BUS_DATA_WIDTH-1 downto 0);
    l_sum_base_price_bus_wdat_strobe : out std_logic_vector(L_SUM_BASE_PRICE_BUS_DATA_WIDTH/8-1 downto 0);
    l_sum_base_price_bus_wdat_last   : out std_logic;
    l_sum_base_price_cmd_valid       : in  std_logic;
    l_sum_base_price_cmd_ready       : out std_logic;
    l_sum_base_price_cmd_firstIdx    : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_sum_base_price_cmd_lastIdx     : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_sum_base_price_cmd_ctrl        : in  std_logic_vector(L_SUM_BASE_PRICE_BUS_ADDR_WIDTH-1 downto 0);
    l_sum_base_price_cmd_tag         : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_sum_base_price_unl_valid       : out std_logic;
    l_sum_base_price_unl_ready       : in  std_logic;
    l_sum_base_price_unl_tag         : out std_logic_vector(TAG_WIDTH-1 downto 0);
    l_sum_disc_price_valid           : in  std_logic;
    l_sum_disc_price_ready           : out std_logic;
    l_sum_disc_price_dvalid          : in  std_logic;
    l_sum_disc_price_last            : in  std_logic;
    l_sum_disc_price                 : in  std_logic_vector(63 downto 0);
    l_sum_disc_price_bus_wreq_valid  : out std_logic;
    l_sum_disc_price_bus_wreq_ready  : in  std_logic;
    l_sum_disc_price_bus_wreq_addr   : out std_logic_vector(L_SUM_DISC_PRICE_BUS_ADDR_WIDTH-1 downto 0);
    l_sum_disc_price_bus_wreq_len    : out std_logic_vector(L_SUM_DISC_PRICE_BUS_LEN_WIDTH-1 downto 0);
    l_sum_disc_price_bus_wdat_valid  : out std_logic;
    l_sum_disc_price_bus_wdat_ready  : in  std_logic;
    l_sum_disc_price_bus_wdat_data   : out std_logic_vector(L_SUM_DISC_PRICE_BUS_DATA_WIDTH-1 downto 0);
    l_sum_disc_price_bus_wdat_strobe : out std_logic_vector(L_SUM_DISC_PRICE_BUS_DATA_WIDTH/8-1 downto 0);
    l_sum_disc_price_bus_wdat_last   : out std_logic;
    l_sum_disc_price_cmd_valid       : in  std_logic;
    l_sum_disc_price_cmd_ready       : out std_logic;
    l_sum_disc_price_cmd_firstIdx    : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_sum_disc_price_cmd_lastIdx     : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_sum_disc_price_cmd_ctrl        : in  std_logic_vector(L_SUM_DISC_PRICE_BUS_ADDR_WIDTH-1 downto 0);
    l_sum_disc_price_cmd_tag         : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_sum_disc_price_unl_valid       : out std_logic;
    l_sum_disc_price_unl_ready       : in  std_logic;
    l_sum_disc_price_unl_tag         : out std_logic_vector(TAG_WIDTH-1 downto 0);
    l_sum_charge_valid               : in  std_logic;
    l_sum_charge_ready               : out std_logic;
    l_sum_charge_dvalid              : in  std_logic;
    l_sum_charge_last                : in  std_logic;
    l_sum_charge                     : in  std_logic_vector(63 downto 0);
    l_sum_charge_bus_wreq_valid      : out std_logic;
    l_sum_charge_bus_wreq_ready      : in  std_logic;
    l_sum_charge_bus_wreq_addr       : out std_logic_vector(L_SUM_CHARGE_BUS_ADDR_WIDTH-1 downto 0);
    l_sum_charge_bus_wreq_len        : out std_logic_vector(L_SUM_CHARGE_BUS_LEN_WIDTH-1 downto 0);
    l_sum_charge_bus_wdat_valid      : out std_logic;
    l_sum_charge_bus_wdat_ready      : in  std_logic;
    l_sum_charge_bus_wdat_data       : out std_logic_vector(L_SUM_CHARGE_BUS_DATA_WIDTH-1 downto 0);
    l_sum_charge_bus_wdat_strobe     : out std_logic_vector(L_SUM_CHARGE_BUS_DATA_WIDTH/8-1 downto 0);
    l_sum_charge_bus_wdat_last       : out std_logic;
    l_sum_charge_cmd_valid           : in  std_logic;
    l_sum_charge_cmd_ready           : out std_logic;
    l_sum_charge_cmd_firstIdx        : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_sum_charge_cmd_lastIdx         : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_sum_charge_cmd_ctrl            : in  std_logic_vector(L_SUM_CHARGE_BUS_ADDR_WIDTH-1 downto 0);
    l_sum_charge_cmd_tag             : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_sum_charge_unl_valid           : out std_logic;
    l_sum_charge_unl_ready           : in  std_logic;
    l_sum_charge_unl_tag             : out std_logic_vector(TAG_WIDTH-1 downto 0);
    l_avg_qty_valid                  : in  std_logic;
    l_avg_qty_ready                  : out std_logic;
    l_avg_qty_dvalid                 : in  std_logic;
    l_avg_qty_last                   : in  std_logic;
    l_avg_qty                        : in  std_logic_vector(63 downto 0);
    l_avg_qty_bus_wreq_valid         : out std_logic;
    l_avg_qty_bus_wreq_ready         : in  std_logic;
    l_avg_qty_bus_wreq_addr          : out std_logic_vector(L_AVG_QTY_BUS_ADDR_WIDTH-1 downto 0);
    l_avg_qty_bus_wreq_len           : out std_logic_vector(L_AVG_QTY_BUS_LEN_WIDTH-1 downto 0);
    l_avg_qty_bus_wdat_valid         : out std_logic;
    l_avg_qty_bus_wdat_ready         : in  std_logic;
    l_avg_qty_bus_wdat_data          : out std_logic_vector(L_AVG_QTY_BUS_DATA_WIDTH-1 downto 0);
    l_avg_qty_bus_wdat_strobe        : out std_logic_vector(L_AVG_QTY_BUS_DATA_WIDTH/8-1 downto 0);
    l_avg_qty_bus_wdat_last          : out std_logic;
    l_avg_qty_cmd_valid              : in  std_logic;
    l_avg_qty_cmd_ready              : out std_logic;
    l_avg_qty_cmd_firstIdx           : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_avg_qty_cmd_lastIdx            : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_avg_qty_cmd_ctrl               : in  std_logic_vector(L_AVG_QTY_BUS_ADDR_WIDTH-1 downto 0);
    l_avg_qty_cmd_tag                : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_avg_qty_unl_valid              : out std_logic;
    l_avg_qty_unl_ready              : in  std_logic;
    l_avg_qty_unl_tag                : out std_logic_vector(TAG_WIDTH-1 downto 0);
    l_avg_price_valid                : in  std_logic;
    l_avg_price_ready                : out std_logic;
    l_avg_price_dvalid               : in  std_logic;
    l_avg_price_last                 : in  std_logic;
    l_avg_price                      : in  std_logic_vector(63 downto 0);
    l_avg_price_bus_wreq_valid       : out std_logic;
    l_avg_price_bus_wreq_ready       : in  std_logic;
    l_avg_price_bus_wreq_addr        : out std_logic_vector(L_AVG_PRICE_BUS_ADDR_WIDTH-1 downto 0);
    l_avg_price_bus_wreq_len         : out std_logic_vector(L_AVG_PRICE_BUS_LEN_WIDTH-1 downto 0);
    l_avg_price_bus_wdat_valid       : out std_logic;
    l_avg_price_bus_wdat_ready       : in  std_logic;
    l_avg_price_bus_wdat_data        : out std_logic_vector(L_AVG_PRICE_BUS_DATA_WIDTH-1 downto 0);
    l_avg_price_bus_wdat_strobe      : out std_logic_vector(L_AVG_PRICE_BUS_DATA_WIDTH/8-1 downto 0);
    l_avg_price_bus_wdat_last        : out std_logic;
    l_avg_price_cmd_valid            : in  std_logic;
    l_avg_price_cmd_ready            : out std_logic;
    l_avg_price_cmd_firstIdx         : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_avg_price_cmd_lastIdx          : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_avg_price_cmd_ctrl             : in  std_logic_vector(L_AVG_PRICE_BUS_ADDR_WIDTH-1 downto 0);
    l_avg_price_cmd_tag              : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_avg_price_unl_valid            : out std_logic;
    l_avg_price_unl_ready            : in  std_logic;
    l_avg_price_unl_tag              : out std_logic_vector(TAG_WIDTH-1 downto 0);
    l_avg_disc_valid                 : in  std_logic;
    l_avg_disc_ready                 : out std_logic;
    l_avg_disc_dvalid                : in  std_logic;
    l_avg_disc_last                  : in  std_logic;
    l_avg_disc                       : in  std_logic_vector(63 downto 0);
    l_avg_disc_bus_wreq_valid        : out std_logic;
    l_avg_disc_bus_wreq_ready        : in  std_logic;
    l_avg_disc_bus_wreq_addr         : out std_logic_vector(L_AVG_DISC_BUS_ADDR_WIDTH-1 downto 0);
    l_avg_disc_bus_wreq_len          : out std_logic_vector(L_AVG_DISC_BUS_LEN_WIDTH-1 downto 0);
    l_avg_disc_bus_wdat_valid        : out std_logic;
    l_avg_disc_bus_wdat_ready        : in  std_logic;
    l_avg_disc_bus_wdat_data         : out std_logic_vector(L_AVG_DISC_BUS_DATA_WIDTH-1 downto 0);
    l_avg_disc_bus_wdat_strobe       : out std_logic_vector(L_AVG_DISC_BUS_DATA_WIDTH/8-1 downto 0);
    l_avg_disc_bus_wdat_last         : out std_logic;
    l_avg_disc_cmd_valid             : in  std_logic;
    l_avg_disc_cmd_ready             : out std_logic;
    l_avg_disc_cmd_firstIdx          : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_avg_disc_cmd_lastIdx           : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_avg_disc_cmd_ctrl              : in  std_logic_vector(L_AVG_DISC_BUS_ADDR_WIDTH-1 downto 0);
    l_avg_disc_cmd_tag               : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_avg_disc_unl_valid             : out std_logic;
    l_avg_disc_unl_ready             : in  std_logic;
    l_avg_disc_unl_tag               : out std_logic_vector(TAG_WIDTH-1 downto 0);
    l_count_order_valid              : in  std_logic;
    l_count_order_ready              : out std_logic;
    l_count_order_dvalid             : in  std_logic;
    l_count_order_last               : in  std_logic;
    l_count_order                    : in  std_logic_vector(63 downto 0);
    l_count_order_bus_wreq_valid     : out std_logic;
    l_count_order_bus_wreq_ready     : in  std_logic;
    l_count_order_bus_wreq_addr      : out std_logic_vector(L_COUNT_ORDER_BUS_ADDR_WIDTH-1 downto 0);
    l_count_order_bus_wreq_len       : out std_logic_vector(L_COUNT_ORDER_BUS_LEN_WIDTH-1 downto 0);
    l_count_order_bus_wdat_valid     : out std_logic;
    l_count_order_bus_wdat_ready     : in  std_logic;
    l_count_order_bus_wdat_data      : out std_logic_vector(L_COUNT_ORDER_BUS_DATA_WIDTH-1 downto 0);
    l_count_order_bus_wdat_strobe    : out std_logic_vector(L_COUNT_ORDER_BUS_DATA_WIDTH/8-1 downto 0);
    l_count_order_bus_wdat_last      : out std_logic;
    l_count_order_cmd_valid          : in  std_logic;
    l_count_order_cmd_ready          : out std_logic;
    l_count_order_cmd_firstIdx       : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_count_order_cmd_lastIdx        : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_count_order_cmd_ctrl           : in  std_logic_vector(L_COUNT_ORDER_BUS_ADDR_WIDTH-1 downto 0);
    l_count_order_cmd_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_count_order_unl_valid          : out std_logic;
    l_count_order_unl_ready          : in  std_logic;
    l_count_order_unl_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0)
  );
end entity;

architecture Implementation of PriceSummaryWriter_l is
  signal returnflag_o_inst_cmd_valid         : std_logic;
  signal returnflag_o_inst_cmd_ready         : std_logic;
  signal returnflag_o_inst_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal returnflag_o_inst_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal returnflag_o_inst_cmd_ctrl          : std_logic_vector(L_RETURNFLAG_O_BUS_ADDR_WIDTH*2-1 downto 0);
  signal returnflag_o_inst_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal returnflag_o_inst_unl_valid         : std_logic;
  signal returnflag_o_inst_unl_ready         : std_logic;
  signal returnflag_o_inst_unl_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal returnflag_o_inst_bus_wreq_valid    : std_logic;
  signal returnflag_o_inst_bus_wreq_ready    : std_logic;
  signal returnflag_o_inst_bus_wreq_addr     : std_logic_vector(L_RETURNFLAG_O_BUS_ADDR_WIDTH-1 downto 0);
  signal returnflag_o_inst_bus_wreq_len      : std_logic_vector(L_RETURNFLAG_O_BUS_LEN_WIDTH-1 downto 0);
  signal returnflag_o_inst_bus_wdat_valid    : std_logic;
  signal returnflag_o_inst_bus_wdat_ready    : std_logic;
  signal returnflag_o_inst_bus_wdat_data     : std_logic_vector(L_RETURNFLAG_O_BUS_DATA_WIDTH-1 downto 0);
  signal returnflag_o_inst_bus_wdat_strobe   : std_logic_vector(L_RETURNFLAG_O_BUS_DATA_WIDTH/8-1 downto 0);
  signal returnflag_o_inst_bus_wdat_last     : std_logic;

  signal returnflag_o_inst_in_valid          : std_logic_vector(1 downto 0);
  signal returnflag_o_inst_in_ready          : std_logic_vector(1 downto 0);
  signal returnflag_o_inst_in_data           : std_logic_vector(41 downto 0);
  signal returnflag_o_inst_in_dvalid         : std_logic_vector(1 downto 0);
  signal returnflag_o_inst_in_last           : std_logic_vector(1 downto 0);

  signal linestatus_o_inst_cmd_valid         : std_logic;
  signal linestatus_o_inst_cmd_ready         : std_logic;
  signal linestatus_o_inst_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal linestatus_o_inst_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal linestatus_o_inst_cmd_ctrl          : std_logic_vector(L_LINESTATUS_O_BUS_ADDR_WIDTH*2-1 downto 0);
  signal linestatus_o_inst_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal linestatus_o_inst_unl_valid         : std_logic;
  signal linestatus_o_inst_unl_ready         : std_logic;
  signal linestatus_o_inst_unl_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal linestatus_o_inst_bus_wreq_valid    : std_logic;
  signal linestatus_o_inst_bus_wreq_ready    : std_logic;
  signal linestatus_o_inst_bus_wreq_addr     : std_logic_vector(L_LINESTATUS_O_BUS_ADDR_WIDTH-1 downto 0);
  signal linestatus_o_inst_bus_wreq_len      : std_logic_vector(L_LINESTATUS_O_BUS_LEN_WIDTH-1 downto 0);
  signal linestatus_o_inst_bus_wdat_valid    : std_logic;
  signal linestatus_o_inst_bus_wdat_ready    : std_logic;
  signal linestatus_o_inst_bus_wdat_data     : std_logic_vector(L_LINESTATUS_O_BUS_DATA_WIDTH-1 downto 0);
  signal linestatus_o_inst_bus_wdat_strobe   : std_logic_vector(L_LINESTATUS_O_BUS_DATA_WIDTH/8-1 downto 0);
  signal linestatus_o_inst_bus_wdat_last     : std_logic;

  signal linestatus_o_inst_in_valid          : std_logic_vector(1 downto 0);
  signal linestatus_o_inst_in_ready          : std_logic_vector(1 downto 0);
  signal linestatus_o_inst_in_data           : std_logic_vector(41 downto 0);
  signal linestatus_o_inst_in_dvalid         : std_logic_vector(1 downto 0);
  signal linestatus_o_inst_in_last           : std_logic_vector(1 downto 0);

  signal sum_qty_inst_cmd_valid              : std_logic;
  signal sum_qty_inst_cmd_ready              : std_logic;
  signal sum_qty_inst_cmd_firstIdx           : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal sum_qty_inst_cmd_lastIdx            : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal sum_qty_inst_cmd_ctrl               : std_logic_vector(L_SUM_QTY_BUS_ADDR_WIDTH-1 downto 0);
  signal sum_qty_inst_cmd_tag                : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal sum_qty_inst_unl_valid              : std_logic;
  signal sum_qty_inst_unl_ready              : std_logic;
  signal sum_qty_inst_unl_tag                : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal sum_qty_inst_bus_wreq_valid         : std_logic;
  signal sum_qty_inst_bus_wreq_ready         : std_logic;
  signal sum_qty_inst_bus_wreq_addr          : std_logic_vector(L_SUM_QTY_BUS_ADDR_WIDTH-1 downto 0);
  signal sum_qty_inst_bus_wreq_len           : std_logic_vector(L_SUM_QTY_BUS_LEN_WIDTH-1 downto 0);
  signal sum_qty_inst_bus_wdat_valid         : std_logic;
  signal sum_qty_inst_bus_wdat_ready         : std_logic;
  signal sum_qty_inst_bus_wdat_data          : std_logic_vector(L_SUM_QTY_BUS_DATA_WIDTH-1 downto 0);
  signal sum_qty_inst_bus_wdat_strobe        : std_logic_vector(L_SUM_QTY_BUS_DATA_WIDTH/8-1 downto 0);
  signal sum_qty_inst_bus_wdat_last          : std_logic;

  signal sum_qty_inst_in_valid               : std_logic_vector(0 downto 0);
  signal sum_qty_inst_in_ready               : std_logic_vector(0 downto 0);
  signal sum_qty_inst_in_data                : std_logic_vector(63 downto 0);
  signal sum_qty_inst_in_dvalid              : std_logic_vector(0 downto 0);
  signal sum_qty_inst_in_last                : std_logic_vector(0 downto 0);

  signal sum_base_price_inst_cmd_valid       : std_logic;
  signal sum_base_price_inst_cmd_ready       : std_logic;
  signal sum_base_price_inst_cmd_firstIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal sum_base_price_inst_cmd_lastIdx     : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal sum_base_price_inst_cmd_ctrl        : std_logic_vector(L_SUM_BASE_PRICE_BUS_ADDR_WIDTH-1 downto 0);
  signal sum_base_price_inst_cmd_tag         : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal sum_base_price_inst_unl_valid       : std_logic;
  signal sum_base_price_inst_unl_ready       : std_logic;
  signal sum_base_price_inst_unl_tag         : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal sum_base_price_inst_bus_wreq_valid  : std_logic;
  signal sum_base_price_inst_bus_wreq_ready  : std_logic;
  signal sum_base_price_inst_bus_wreq_addr   : std_logic_vector(L_SUM_BASE_PRICE_BUS_ADDR_WIDTH-1 downto 0);
  signal sum_base_price_inst_bus_wreq_len    : std_logic_vector(L_SUM_BASE_PRICE_BUS_LEN_WIDTH-1 downto 0);
  signal sum_base_price_inst_bus_wdat_valid  : std_logic;
  signal sum_base_price_inst_bus_wdat_ready  : std_logic;
  signal sum_base_price_inst_bus_wdat_data   : std_logic_vector(L_SUM_BASE_PRICE_BUS_DATA_WIDTH-1 downto 0);
  signal sum_base_price_inst_bus_wdat_strobe : std_logic_vector(L_SUM_BASE_PRICE_BUS_DATA_WIDTH/8-1 downto 0);
  signal sum_base_price_inst_bus_wdat_last   : std_logic;

  signal sum_base_price_inst_in_valid        : std_logic_vector(0 downto 0);
  signal sum_base_price_inst_in_ready        : std_logic_vector(0 downto 0);
  signal sum_base_price_inst_in_data         : std_logic_vector(63 downto 0);
  signal sum_base_price_inst_in_dvalid       : std_logic_vector(0 downto 0);
  signal sum_base_price_inst_in_last         : std_logic_vector(0 downto 0);

  signal sum_disc_price_inst_cmd_valid       : std_logic;
  signal sum_disc_price_inst_cmd_ready       : std_logic;
  signal sum_disc_price_inst_cmd_firstIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal sum_disc_price_inst_cmd_lastIdx     : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal sum_disc_price_inst_cmd_ctrl        : std_logic_vector(L_SUM_DISC_PRICE_BUS_ADDR_WIDTH-1 downto 0);
  signal sum_disc_price_inst_cmd_tag         : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal sum_disc_price_inst_unl_valid       : std_logic;
  signal sum_disc_price_inst_unl_ready       : std_logic;
  signal sum_disc_price_inst_unl_tag         : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal sum_disc_price_inst_bus_wreq_valid  : std_logic;
  signal sum_disc_price_inst_bus_wreq_ready  : std_logic;
  signal sum_disc_price_inst_bus_wreq_addr   : std_logic_vector(L_SUM_DISC_PRICE_BUS_ADDR_WIDTH-1 downto 0);
  signal sum_disc_price_inst_bus_wreq_len    : std_logic_vector(L_SUM_DISC_PRICE_BUS_LEN_WIDTH-1 downto 0);
  signal sum_disc_price_inst_bus_wdat_valid  : std_logic;
  signal sum_disc_price_inst_bus_wdat_ready  : std_logic;
  signal sum_disc_price_inst_bus_wdat_data   : std_logic_vector(L_SUM_DISC_PRICE_BUS_DATA_WIDTH-1 downto 0);
  signal sum_disc_price_inst_bus_wdat_strobe : std_logic_vector(L_SUM_DISC_PRICE_BUS_DATA_WIDTH/8-1 downto 0);
  signal sum_disc_price_inst_bus_wdat_last   : std_logic;

  signal sum_disc_price_inst_in_valid        : std_logic_vector(0 downto 0);
  signal sum_disc_price_inst_in_ready        : std_logic_vector(0 downto 0);
  signal sum_disc_price_inst_in_data         : std_logic_vector(63 downto 0);
  signal sum_disc_price_inst_in_dvalid       : std_logic_vector(0 downto 0);
  signal sum_disc_price_inst_in_last         : std_logic_vector(0 downto 0);

  signal sum_charge_inst_cmd_valid           : std_logic;
  signal sum_charge_inst_cmd_ready           : std_logic;
  signal sum_charge_inst_cmd_firstIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal sum_charge_inst_cmd_lastIdx         : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal sum_charge_inst_cmd_ctrl            : std_logic_vector(L_SUM_CHARGE_BUS_ADDR_WIDTH-1 downto 0);
  signal sum_charge_inst_cmd_tag             : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal sum_charge_inst_unl_valid           : std_logic;
  signal sum_charge_inst_unl_ready           : std_logic;
  signal sum_charge_inst_unl_tag             : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal sum_charge_inst_bus_wreq_valid      : std_logic;
  signal sum_charge_inst_bus_wreq_ready      : std_logic;
  signal sum_charge_inst_bus_wreq_addr       : std_logic_vector(L_SUM_CHARGE_BUS_ADDR_WIDTH-1 downto 0);
  signal sum_charge_inst_bus_wreq_len        : std_logic_vector(L_SUM_CHARGE_BUS_LEN_WIDTH-1 downto 0);
  signal sum_charge_inst_bus_wdat_valid      : std_logic;
  signal sum_charge_inst_bus_wdat_ready      : std_logic;
  signal sum_charge_inst_bus_wdat_data       : std_logic_vector(L_SUM_CHARGE_BUS_DATA_WIDTH-1 downto 0);
  signal sum_charge_inst_bus_wdat_strobe     : std_logic_vector(L_SUM_CHARGE_BUS_DATA_WIDTH/8-1 downto 0);
  signal sum_charge_inst_bus_wdat_last       : std_logic;

  signal sum_charge_inst_in_valid            : std_logic_vector(0 downto 0);
  signal sum_charge_inst_in_ready            : std_logic_vector(0 downto 0);
  signal sum_charge_inst_in_data             : std_logic_vector(63 downto 0);
  signal sum_charge_inst_in_dvalid           : std_logic_vector(0 downto 0);
  signal sum_charge_inst_in_last             : std_logic_vector(0 downto 0);

  signal avg_qty_inst_cmd_valid              : std_logic;
  signal avg_qty_inst_cmd_ready              : std_logic;
  signal avg_qty_inst_cmd_firstIdx           : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal avg_qty_inst_cmd_lastIdx            : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal avg_qty_inst_cmd_ctrl               : std_logic_vector(L_AVG_QTY_BUS_ADDR_WIDTH-1 downto 0);
  signal avg_qty_inst_cmd_tag                : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal avg_qty_inst_unl_valid              : std_logic;
  signal avg_qty_inst_unl_ready              : std_logic;
  signal avg_qty_inst_unl_tag                : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal avg_qty_inst_bus_wreq_valid         : std_logic;
  signal avg_qty_inst_bus_wreq_ready         : std_logic;
  signal avg_qty_inst_bus_wreq_addr          : std_logic_vector(L_AVG_QTY_BUS_ADDR_WIDTH-1 downto 0);
  signal avg_qty_inst_bus_wreq_len           : std_logic_vector(L_AVG_QTY_BUS_LEN_WIDTH-1 downto 0);
  signal avg_qty_inst_bus_wdat_valid         : std_logic;
  signal avg_qty_inst_bus_wdat_ready         : std_logic;
  signal avg_qty_inst_bus_wdat_data          : std_logic_vector(L_AVG_QTY_BUS_DATA_WIDTH-1 downto 0);
  signal avg_qty_inst_bus_wdat_strobe        : std_logic_vector(L_AVG_QTY_BUS_DATA_WIDTH/8-1 downto 0);
  signal avg_qty_inst_bus_wdat_last          : std_logic;

  signal avg_qty_inst_in_valid               : std_logic_vector(0 downto 0);
  signal avg_qty_inst_in_ready               : std_logic_vector(0 downto 0);
  signal avg_qty_inst_in_data                : std_logic_vector(63 downto 0);
  signal avg_qty_inst_in_dvalid              : std_logic_vector(0 downto 0);
  signal avg_qty_inst_in_last                : std_logic_vector(0 downto 0);

  signal avg_price_inst_cmd_valid            : std_logic;
  signal avg_price_inst_cmd_ready            : std_logic;
  signal avg_price_inst_cmd_firstIdx         : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal avg_price_inst_cmd_lastIdx          : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal avg_price_inst_cmd_ctrl             : std_logic_vector(L_AVG_PRICE_BUS_ADDR_WIDTH-1 downto 0);
  signal avg_price_inst_cmd_tag              : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal avg_price_inst_unl_valid            : std_logic;
  signal avg_price_inst_unl_ready            : std_logic;
  signal avg_price_inst_unl_tag              : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal avg_price_inst_bus_wreq_valid       : std_logic;
  signal avg_price_inst_bus_wreq_ready       : std_logic;
  signal avg_price_inst_bus_wreq_addr        : std_logic_vector(L_AVG_PRICE_BUS_ADDR_WIDTH-1 downto 0);
  signal avg_price_inst_bus_wreq_len         : std_logic_vector(L_AVG_PRICE_BUS_LEN_WIDTH-1 downto 0);
  signal avg_price_inst_bus_wdat_valid       : std_logic;
  signal avg_price_inst_bus_wdat_ready       : std_logic;
  signal avg_price_inst_bus_wdat_data        : std_logic_vector(L_AVG_PRICE_BUS_DATA_WIDTH-1 downto 0);
  signal avg_price_inst_bus_wdat_strobe      : std_logic_vector(L_AVG_PRICE_BUS_DATA_WIDTH/8-1 downto 0);
  signal avg_price_inst_bus_wdat_last        : std_logic;

  signal avg_price_inst_in_valid             : std_logic_vector(0 downto 0);
  signal avg_price_inst_in_ready             : std_logic_vector(0 downto 0);
  signal avg_price_inst_in_data              : std_logic_vector(63 downto 0);
  signal avg_price_inst_in_dvalid            : std_logic_vector(0 downto 0);
  signal avg_price_inst_in_last              : std_logic_vector(0 downto 0);

  signal avg_disc_inst_cmd_valid             : std_logic;
  signal avg_disc_inst_cmd_ready             : std_logic;
  signal avg_disc_inst_cmd_firstIdx          : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal avg_disc_inst_cmd_lastIdx           : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal avg_disc_inst_cmd_ctrl              : std_logic_vector(L_AVG_DISC_BUS_ADDR_WIDTH-1 downto 0);
  signal avg_disc_inst_cmd_tag               : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal avg_disc_inst_unl_valid             : std_logic;
  signal avg_disc_inst_unl_ready             : std_logic;
  signal avg_disc_inst_unl_tag               : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal avg_disc_inst_bus_wreq_valid        : std_logic;
  signal avg_disc_inst_bus_wreq_ready        : std_logic;
  signal avg_disc_inst_bus_wreq_addr         : std_logic_vector(L_AVG_DISC_BUS_ADDR_WIDTH-1 downto 0);
  signal avg_disc_inst_bus_wreq_len          : std_logic_vector(L_AVG_DISC_BUS_LEN_WIDTH-1 downto 0);
  signal avg_disc_inst_bus_wdat_valid        : std_logic;
  signal avg_disc_inst_bus_wdat_ready        : std_logic;
  signal avg_disc_inst_bus_wdat_data         : std_logic_vector(L_AVG_DISC_BUS_DATA_WIDTH-1 downto 0);
  signal avg_disc_inst_bus_wdat_strobe       : std_logic_vector(L_AVG_DISC_BUS_DATA_WIDTH/8-1 downto 0);
  signal avg_disc_inst_bus_wdat_last         : std_logic;

  signal avg_disc_inst_in_valid              : std_logic_vector(0 downto 0);
  signal avg_disc_inst_in_ready              : std_logic_vector(0 downto 0);
  signal avg_disc_inst_in_data               : std_logic_vector(63 downto 0);
  signal avg_disc_inst_in_dvalid             : std_logic_vector(0 downto 0);
  signal avg_disc_inst_in_last               : std_logic_vector(0 downto 0);

  signal count_order_inst_cmd_valid          : std_logic;
  signal count_order_inst_cmd_ready          : std_logic;
  signal count_order_inst_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal count_order_inst_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal count_order_inst_cmd_ctrl           : std_logic_vector(L_COUNT_ORDER_BUS_ADDR_WIDTH-1 downto 0);
  signal count_order_inst_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal count_order_inst_unl_valid          : std_logic;
  signal count_order_inst_unl_ready          : std_logic;
  signal count_order_inst_unl_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal count_order_inst_bus_wreq_valid     : std_logic;
  signal count_order_inst_bus_wreq_ready     : std_logic;
  signal count_order_inst_bus_wreq_addr      : std_logic_vector(L_COUNT_ORDER_BUS_ADDR_WIDTH-1 downto 0);
  signal count_order_inst_bus_wreq_len       : std_logic_vector(L_COUNT_ORDER_BUS_LEN_WIDTH-1 downto 0);
  signal count_order_inst_bus_wdat_valid     : std_logic;
  signal count_order_inst_bus_wdat_ready     : std_logic;
  signal count_order_inst_bus_wdat_data      : std_logic_vector(L_COUNT_ORDER_BUS_DATA_WIDTH-1 downto 0);
  signal count_order_inst_bus_wdat_strobe    : std_logic_vector(L_COUNT_ORDER_BUS_DATA_WIDTH/8-1 downto 0);
  signal count_order_inst_bus_wdat_last      : std_logic;

  signal count_order_inst_in_valid           : std_logic_vector(0 downto 0);
  signal count_order_inst_in_ready           : std_logic_vector(0 downto 0);
  signal count_order_inst_in_data            : std_logic_vector(63 downto 0);
  signal count_order_inst_in_dvalid          : std_logic_vector(0 downto 0);
  signal count_order_inst_in_last            : std_logic_vector(0 downto 0);

begin
  returnflag_o_inst : ArrayWriter
    generic map (
      BUS_ADDR_WIDTH     => L_RETURNFLAG_O_BUS_ADDR_WIDTH,
      BUS_DATA_WIDTH     => L_RETURNFLAG_O_BUS_DATA_WIDTH,
      BUS_LEN_WIDTH      => L_RETURNFLAG_O_BUS_LEN_WIDTH,
      BUS_BURST_STEP_LEN => L_RETURNFLAG_O_BUS_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN  => L_RETURNFLAG_O_BUS_BURST_MAX_LEN,
      INDEX_WIDTH        => INDEX_WIDTH,
      CFG                => "listprim(8)",
      CMD_TAG_ENABLE     => true,
      CMD_TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      bcd_clk         => bcd_clk,
      bcd_reset       => bcd_reset,
      kcd_clk         => kcd_clk,
      kcd_reset       => kcd_reset,
      cmd_valid       => returnflag_o_inst_cmd_valid,
      cmd_ready       => returnflag_o_inst_cmd_ready,
      cmd_firstIdx    => returnflag_o_inst_cmd_firstIdx,
      cmd_lastIdx     => returnflag_o_inst_cmd_lastIdx,
      cmd_ctrl        => returnflag_o_inst_cmd_ctrl,
      cmd_tag         => returnflag_o_inst_cmd_tag,
      unl_valid       => returnflag_o_inst_unl_valid,
      unl_ready       => returnflag_o_inst_unl_ready,
      unl_tag         => returnflag_o_inst_unl_tag,
      bus_wreq_valid  => returnflag_o_inst_bus_wreq_valid,
      bus_wreq_ready  => returnflag_o_inst_bus_wreq_ready,
      bus_wreq_addr   => returnflag_o_inst_bus_wreq_addr,
      bus_wreq_len    => returnflag_o_inst_bus_wreq_len,
      bus_wdat_valid  => returnflag_o_inst_bus_wdat_valid,
      bus_wdat_ready  => returnflag_o_inst_bus_wdat_ready,
      bus_wdat_data   => returnflag_o_inst_bus_wdat_data,
      bus_wdat_strobe => returnflag_o_inst_bus_wdat_strobe,
      bus_wdat_last   => returnflag_o_inst_bus_wdat_last,
      in_valid        => returnflag_o_inst_in_valid,
      in_ready        => returnflag_o_inst_in_ready,
      in_data         => returnflag_o_inst_in_data,
      in_dvalid       => returnflag_o_inst_in_dvalid,
      in_last         => returnflag_o_inst_in_last
    );

  linestatus_o_inst : ArrayWriter
    generic map (
      BUS_ADDR_WIDTH     => L_LINESTATUS_O_BUS_ADDR_WIDTH,
      BUS_DATA_WIDTH     => L_LINESTATUS_O_BUS_DATA_WIDTH,
      BUS_LEN_WIDTH      => L_LINESTATUS_O_BUS_LEN_WIDTH,
      BUS_BURST_STEP_LEN => L_LINESTATUS_O_BUS_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN  => L_LINESTATUS_O_BUS_BURST_MAX_LEN,
      INDEX_WIDTH        => INDEX_WIDTH,
      CFG                => "listprim(8)",
      CMD_TAG_ENABLE     => true,
      CMD_TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      bcd_clk         => bcd_clk,
      bcd_reset       => bcd_reset,
      kcd_clk         => kcd_clk,
      kcd_reset       => kcd_reset,
      cmd_valid       => linestatus_o_inst_cmd_valid,
      cmd_ready       => linestatus_o_inst_cmd_ready,
      cmd_firstIdx    => linestatus_o_inst_cmd_firstIdx,
      cmd_lastIdx     => linestatus_o_inst_cmd_lastIdx,
      cmd_ctrl        => linestatus_o_inst_cmd_ctrl,
      cmd_tag         => linestatus_o_inst_cmd_tag,
      unl_valid       => linestatus_o_inst_unl_valid,
      unl_ready       => linestatus_o_inst_unl_ready,
      unl_tag         => linestatus_o_inst_unl_tag,
      bus_wreq_valid  => linestatus_o_inst_bus_wreq_valid,
      bus_wreq_ready  => linestatus_o_inst_bus_wreq_ready,
      bus_wreq_addr   => linestatus_o_inst_bus_wreq_addr,
      bus_wreq_len    => linestatus_o_inst_bus_wreq_len,
      bus_wdat_valid  => linestatus_o_inst_bus_wdat_valid,
      bus_wdat_ready  => linestatus_o_inst_bus_wdat_ready,
      bus_wdat_data   => linestatus_o_inst_bus_wdat_data,
      bus_wdat_strobe => linestatus_o_inst_bus_wdat_strobe,
      bus_wdat_last   => linestatus_o_inst_bus_wdat_last,
      in_valid        => linestatus_o_inst_in_valid,
      in_ready        => linestatus_o_inst_in_ready,
      in_data         => linestatus_o_inst_in_data,
      in_dvalid       => linestatus_o_inst_in_dvalid,
      in_last         => linestatus_o_inst_in_last
    );

  sum_qty_inst : ArrayWriter
    generic map (
      BUS_ADDR_WIDTH     => L_SUM_QTY_BUS_ADDR_WIDTH,
      BUS_DATA_WIDTH     => L_SUM_QTY_BUS_DATA_WIDTH,
      BUS_LEN_WIDTH      => L_SUM_QTY_BUS_LEN_WIDTH,
      BUS_BURST_STEP_LEN => L_SUM_QTY_BUS_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN  => L_SUM_QTY_BUS_BURST_MAX_LEN,
      INDEX_WIDTH        => INDEX_WIDTH,
      CFG                => "prim(64)",
      CMD_TAG_ENABLE     => true,
      CMD_TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      bcd_clk         => bcd_clk,
      bcd_reset       => bcd_reset,
      kcd_clk         => kcd_clk,
      kcd_reset       => kcd_reset,
      cmd_valid       => sum_qty_inst_cmd_valid,
      cmd_ready       => sum_qty_inst_cmd_ready,
      cmd_firstIdx    => sum_qty_inst_cmd_firstIdx,
      cmd_lastIdx     => sum_qty_inst_cmd_lastIdx,
      cmd_ctrl        => sum_qty_inst_cmd_ctrl,
      cmd_tag         => sum_qty_inst_cmd_tag,
      unl_valid       => sum_qty_inst_unl_valid,
      unl_ready       => sum_qty_inst_unl_ready,
      unl_tag         => sum_qty_inst_unl_tag,
      bus_wreq_valid  => sum_qty_inst_bus_wreq_valid,
      bus_wreq_ready  => sum_qty_inst_bus_wreq_ready,
      bus_wreq_addr   => sum_qty_inst_bus_wreq_addr,
      bus_wreq_len    => sum_qty_inst_bus_wreq_len,
      bus_wdat_valid  => sum_qty_inst_bus_wdat_valid,
      bus_wdat_ready  => sum_qty_inst_bus_wdat_ready,
      bus_wdat_data   => sum_qty_inst_bus_wdat_data,
      bus_wdat_strobe => sum_qty_inst_bus_wdat_strobe,
      bus_wdat_last   => sum_qty_inst_bus_wdat_last,
      in_valid        => sum_qty_inst_in_valid,
      in_ready        => sum_qty_inst_in_ready,
      in_data         => sum_qty_inst_in_data,
      in_dvalid       => sum_qty_inst_in_dvalid,
      in_last         => sum_qty_inst_in_last
    );

  sum_base_price_inst : ArrayWriter
    generic map (
      BUS_ADDR_WIDTH     => L_SUM_BASE_PRICE_BUS_ADDR_WIDTH,
      BUS_DATA_WIDTH     => L_SUM_BASE_PRICE_BUS_DATA_WIDTH,
      BUS_LEN_WIDTH      => L_SUM_BASE_PRICE_BUS_LEN_WIDTH,
      BUS_BURST_STEP_LEN => L_SUM_BASE_PRICE_BUS_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN  => L_SUM_BASE_PRICE_BUS_BURST_MAX_LEN,
      INDEX_WIDTH        => INDEX_WIDTH,
      CFG                => "prim(64)",
      CMD_TAG_ENABLE     => true,
      CMD_TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      bcd_clk         => bcd_clk,
      bcd_reset       => bcd_reset,
      kcd_clk         => kcd_clk,
      kcd_reset       => kcd_reset,
      cmd_valid       => sum_base_price_inst_cmd_valid,
      cmd_ready       => sum_base_price_inst_cmd_ready,
      cmd_firstIdx    => sum_base_price_inst_cmd_firstIdx,
      cmd_lastIdx     => sum_base_price_inst_cmd_lastIdx,
      cmd_ctrl        => sum_base_price_inst_cmd_ctrl,
      cmd_tag         => sum_base_price_inst_cmd_tag,
      unl_valid       => sum_base_price_inst_unl_valid,
      unl_ready       => sum_base_price_inst_unl_ready,
      unl_tag         => sum_base_price_inst_unl_tag,
      bus_wreq_valid  => sum_base_price_inst_bus_wreq_valid,
      bus_wreq_ready  => sum_base_price_inst_bus_wreq_ready,
      bus_wreq_addr   => sum_base_price_inst_bus_wreq_addr,
      bus_wreq_len    => sum_base_price_inst_bus_wreq_len,
      bus_wdat_valid  => sum_base_price_inst_bus_wdat_valid,
      bus_wdat_ready  => sum_base_price_inst_bus_wdat_ready,
      bus_wdat_data   => sum_base_price_inst_bus_wdat_data,
      bus_wdat_strobe => sum_base_price_inst_bus_wdat_strobe,
      bus_wdat_last   => sum_base_price_inst_bus_wdat_last,
      in_valid        => sum_base_price_inst_in_valid,
      in_ready        => sum_base_price_inst_in_ready,
      in_data         => sum_base_price_inst_in_data,
      in_dvalid       => sum_base_price_inst_in_dvalid,
      in_last         => sum_base_price_inst_in_last
    );

  sum_disc_price_inst : ArrayWriter
    generic map (
      BUS_ADDR_WIDTH     => L_SUM_DISC_PRICE_BUS_ADDR_WIDTH,
      BUS_DATA_WIDTH     => L_SUM_DISC_PRICE_BUS_DATA_WIDTH,
      BUS_LEN_WIDTH      => L_SUM_DISC_PRICE_BUS_LEN_WIDTH,
      BUS_BURST_STEP_LEN => L_SUM_DISC_PRICE_BUS_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN  => L_SUM_DISC_PRICE_BUS_BURST_MAX_LEN,
      INDEX_WIDTH        => INDEX_WIDTH,
      CFG                => "prim(64)",
      CMD_TAG_ENABLE     => true,
      CMD_TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      bcd_clk         => bcd_clk,
      bcd_reset       => bcd_reset,
      kcd_clk         => kcd_clk,
      kcd_reset       => kcd_reset,
      cmd_valid       => sum_disc_price_inst_cmd_valid,
      cmd_ready       => sum_disc_price_inst_cmd_ready,
      cmd_firstIdx    => sum_disc_price_inst_cmd_firstIdx,
      cmd_lastIdx     => sum_disc_price_inst_cmd_lastIdx,
      cmd_ctrl        => sum_disc_price_inst_cmd_ctrl,
      cmd_tag         => sum_disc_price_inst_cmd_tag,
      unl_valid       => sum_disc_price_inst_unl_valid,
      unl_ready       => sum_disc_price_inst_unl_ready,
      unl_tag         => sum_disc_price_inst_unl_tag,
      bus_wreq_valid  => sum_disc_price_inst_bus_wreq_valid,
      bus_wreq_ready  => sum_disc_price_inst_bus_wreq_ready,
      bus_wreq_addr   => sum_disc_price_inst_bus_wreq_addr,
      bus_wreq_len    => sum_disc_price_inst_bus_wreq_len,
      bus_wdat_valid  => sum_disc_price_inst_bus_wdat_valid,
      bus_wdat_ready  => sum_disc_price_inst_bus_wdat_ready,
      bus_wdat_data   => sum_disc_price_inst_bus_wdat_data,
      bus_wdat_strobe => sum_disc_price_inst_bus_wdat_strobe,
      bus_wdat_last   => sum_disc_price_inst_bus_wdat_last,
      in_valid        => sum_disc_price_inst_in_valid,
      in_ready        => sum_disc_price_inst_in_ready,
      in_data         => sum_disc_price_inst_in_data,
      in_dvalid       => sum_disc_price_inst_in_dvalid,
      in_last         => sum_disc_price_inst_in_last
    );

  sum_charge_inst : ArrayWriter
    generic map (
      BUS_ADDR_WIDTH     => L_SUM_CHARGE_BUS_ADDR_WIDTH,
      BUS_DATA_WIDTH     => L_SUM_CHARGE_BUS_DATA_WIDTH,
      BUS_LEN_WIDTH      => L_SUM_CHARGE_BUS_LEN_WIDTH,
      BUS_BURST_STEP_LEN => L_SUM_CHARGE_BUS_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN  => L_SUM_CHARGE_BUS_BURST_MAX_LEN,
      INDEX_WIDTH        => INDEX_WIDTH,
      CFG                => "prim(64)",
      CMD_TAG_ENABLE     => true,
      CMD_TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      bcd_clk         => bcd_clk,
      bcd_reset       => bcd_reset,
      kcd_clk         => kcd_clk,
      kcd_reset       => kcd_reset,
      cmd_valid       => sum_charge_inst_cmd_valid,
      cmd_ready       => sum_charge_inst_cmd_ready,
      cmd_firstIdx    => sum_charge_inst_cmd_firstIdx,
      cmd_lastIdx     => sum_charge_inst_cmd_lastIdx,
      cmd_ctrl        => sum_charge_inst_cmd_ctrl,
      cmd_tag         => sum_charge_inst_cmd_tag,
      unl_valid       => sum_charge_inst_unl_valid,
      unl_ready       => sum_charge_inst_unl_ready,
      unl_tag         => sum_charge_inst_unl_tag,
      bus_wreq_valid  => sum_charge_inst_bus_wreq_valid,
      bus_wreq_ready  => sum_charge_inst_bus_wreq_ready,
      bus_wreq_addr   => sum_charge_inst_bus_wreq_addr,
      bus_wreq_len    => sum_charge_inst_bus_wreq_len,
      bus_wdat_valid  => sum_charge_inst_bus_wdat_valid,
      bus_wdat_ready  => sum_charge_inst_bus_wdat_ready,
      bus_wdat_data   => sum_charge_inst_bus_wdat_data,
      bus_wdat_strobe => sum_charge_inst_bus_wdat_strobe,
      bus_wdat_last   => sum_charge_inst_bus_wdat_last,
      in_valid        => sum_charge_inst_in_valid,
      in_ready        => sum_charge_inst_in_ready,
      in_data         => sum_charge_inst_in_data,
      in_dvalid       => sum_charge_inst_in_dvalid,
      in_last         => sum_charge_inst_in_last
    );

  avg_qty_inst : ArrayWriter
    generic map (
      BUS_ADDR_WIDTH     => L_AVG_QTY_BUS_ADDR_WIDTH,
      BUS_DATA_WIDTH     => L_AVG_QTY_BUS_DATA_WIDTH,
      BUS_LEN_WIDTH      => L_AVG_QTY_BUS_LEN_WIDTH,
      BUS_BURST_STEP_LEN => L_AVG_QTY_BUS_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN  => L_AVG_QTY_BUS_BURST_MAX_LEN,
      INDEX_WIDTH        => INDEX_WIDTH,
      CFG                => "prim(64)",
      CMD_TAG_ENABLE     => true,
      CMD_TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      bcd_clk         => bcd_clk,
      bcd_reset       => bcd_reset,
      kcd_clk         => kcd_clk,
      kcd_reset       => kcd_reset,
      cmd_valid       => avg_qty_inst_cmd_valid,
      cmd_ready       => avg_qty_inst_cmd_ready,
      cmd_firstIdx    => avg_qty_inst_cmd_firstIdx,
      cmd_lastIdx     => avg_qty_inst_cmd_lastIdx,
      cmd_ctrl        => avg_qty_inst_cmd_ctrl,
      cmd_tag         => avg_qty_inst_cmd_tag,
      unl_valid       => avg_qty_inst_unl_valid,
      unl_ready       => avg_qty_inst_unl_ready,
      unl_tag         => avg_qty_inst_unl_tag,
      bus_wreq_valid  => avg_qty_inst_bus_wreq_valid,
      bus_wreq_ready  => avg_qty_inst_bus_wreq_ready,
      bus_wreq_addr   => avg_qty_inst_bus_wreq_addr,
      bus_wreq_len    => avg_qty_inst_bus_wreq_len,
      bus_wdat_valid  => avg_qty_inst_bus_wdat_valid,
      bus_wdat_ready  => avg_qty_inst_bus_wdat_ready,
      bus_wdat_data   => avg_qty_inst_bus_wdat_data,
      bus_wdat_strobe => avg_qty_inst_bus_wdat_strobe,
      bus_wdat_last   => avg_qty_inst_bus_wdat_last,
      in_valid        => avg_qty_inst_in_valid,
      in_ready        => avg_qty_inst_in_ready,
      in_data         => avg_qty_inst_in_data,
      in_dvalid       => avg_qty_inst_in_dvalid,
      in_last         => avg_qty_inst_in_last
    );

  avg_price_inst : ArrayWriter
    generic map (
      BUS_ADDR_WIDTH     => L_AVG_PRICE_BUS_ADDR_WIDTH,
      BUS_DATA_WIDTH     => L_AVG_PRICE_BUS_DATA_WIDTH,
      BUS_LEN_WIDTH      => L_AVG_PRICE_BUS_LEN_WIDTH,
      BUS_BURST_STEP_LEN => L_AVG_PRICE_BUS_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN  => L_AVG_PRICE_BUS_BURST_MAX_LEN,
      INDEX_WIDTH        => INDEX_WIDTH,
      CFG                => "prim(64)",
      CMD_TAG_ENABLE     => true,
      CMD_TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      bcd_clk         => bcd_clk,
      bcd_reset       => bcd_reset,
      kcd_clk         => kcd_clk,
      kcd_reset       => kcd_reset,
      cmd_valid       => avg_price_inst_cmd_valid,
      cmd_ready       => avg_price_inst_cmd_ready,
      cmd_firstIdx    => avg_price_inst_cmd_firstIdx,
      cmd_lastIdx     => avg_price_inst_cmd_lastIdx,
      cmd_ctrl        => avg_price_inst_cmd_ctrl,
      cmd_tag         => avg_price_inst_cmd_tag,
      unl_valid       => avg_price_inst_unl_valid,
      unl_ready       => avg_price_inst_unl_ready,
      unl_tag         => avg_price_inst_unl_tag,
      bus_wreq_valid  => avg_price_inst_bus_wreq_valid,
      bus_wreq_ready  => avg_price_inst_bus_wreq_ready,
      bus_wreq_addr   => avg_price_inst_bus_wreq_addr,
      bus_wreq_len    => avg_price_inst_bus_wreq_len,
      bus_wdat_valid  => avg_price_inst_bus_wdat_valid,
      bus_wdat_ready  => avg_price_inst_bus_wdat_ready,
      bus_wdat_data   => avg_price_inst_bus_wdat_data,
      bus_wdat_strobe => avg_price_inst_bus_wdat_strobe,
      bus_wdat_last   => avg_price_inst_bus_wdat_last,
      in_valid        => avg_price_inst_in_valid,
      in_ready        => avg_price_inst_in_ready,
      in_data         => avg_price_inst_in_data,
      in_dvalid       => avg_price_inst_in_dvalid,
      in_last         => avg_price_inst_in_last
    );

  avg_disc_inst : ArrayWriter
    generic map (
      BUS_ADDR_WIDTH     => L_AVG_DISC_BUS_ADDR_WIDTH,
      BUS_DATA_WIDTH     => L_AVG_DISC_BUS_DATA_WIDTH,
      BUS_LEN_WIDTH      => L_AVG_DISC_BUS_LEN_WIDTH,
      BUS_BURST_STEP_LEN => L_AVG_DISC_BUS_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN  => L_AVG_DISC_BUS_BURST_MAX_LEN,
      INDEX_WIDTH        => INDEX_WIDTH,
      CFG                => "prim(64)",
      CMD_TAG_ENABLE     => true,
      CMD_TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      bcd_clk         => bcd_clk,
      bcd_reset       => bcd_reset,
      kcd_clk         => kcd_clk,
      kcd_reset       => kcd_reset,
      cmd_valid       => avg_disc_inst_cmd_valid,
      cmd_ready       => avg_disc_inst_cmd_ready,
      cmd_firstIdx    => avg_disc_inst_cmd_firstIdx,
      cmd_lastIdx     => avg_disc_inst_cmd_lastIdx,
      cmd_ctrl        => avg_disc_inst_cmd_ctrl,
      cmd_tag         => avg_disc_inst_cmd_tag,
      unl_valid       => avg_disc_inst_unl_valid,
      unl_ready       => avg_disc_inst_unl_ready,
      unl_tag         => avg_disc_inst_unl_tag,
      bus_wreq_valid  => avg_disc_inst_bus_wreq_valid,
      bus_wreq_ready  => avg_disc_inst_bus_wreq_ready,
      bus_wreq_addr   => avg_disc_inst_bus_wreq_addr,
      bus_wreq_len    => avg_disc_inst_bus_wreq_len,
      bus_wdat_valid  => avg_disc_inst_bus_wdat_valid,
      bus_wdat_ready  => avg_disc_inst_bus_wdat_ready,
      bus_wdat_data   => avg_disc_inst_bus_wdat_data,
      bus_wdat_strobe => avg_disc_inst_bus_wdat_strobe,
      bus_wdat_last   => avg_disc_inst_bus_wdat_last,
      in_valid        => avg_disc_inst_in_valid,
      in_ready        => avg_disc_inst_in_ready,
      in_data         => avg_disc_inst_in_data,
      in_dvalid       => avg_disc_inst_in_dvalid,
      in_last         => avg_disc_inst_in_last
    );

  count_order_inst : ArrayWriter
    generic map (
      BUS_ADDR_WIDTH     => L_COUNT_ORDER_BUS_ADDR_WIDTH,
      BUS_DATA_WIDTH     => L_COUNT_ORDER_BUS_DATA_WIDTH,
      BUS_LEN_WIDTH      => L_COUNT_ORDER_BUS_LEN_WIDTH,
      BUS_BURST_STEP_LEN => L_COUNT_ORDER_BUS_BURST_STEP_LEN,
      BUS_BURST_MAX_LEN  => L_COUNT_ORDER_BUS_BURST_MAX_LEN,
      INDEX_WIDTH        => INDEX_WIDTH,
      CFG                => "prim(64)",
      CMD_TAG_ENABLE     => true,
      CMD_TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      bcd_clk         => bcd_clk,
      bcd_reset       => bcd_reset,
      kcd_clk         => kcd_clk,
      kcd_reset       => kcd_reset,
      cmd_valid       => count_order_inst_cmd_valid,
      cmd_ready       => count_order_inst_cmd_ready,
      cmd_firstIdx    => count_order_inst_cmd_firstIdx,
      cmd_lastIdx     => count_order_inst_cmd_lastIdx,
      cmd_ctrl        => count_order_inst_cmd_ctrl,
      cmd_tag         => count_order_inst_cmd_tag,
      unl_valid       => count_order_inst_unl_valid,
      unl_ready       => count_order_inst_unl_ready,
      unl_tag         => count_order_inst_unl_tag,
      bus_wreq_valid  => count_order_inst_bus_wreq_valid,
      bus_wreq_ready  => count_order_inst_bus_wreq_ready,
      bus_wreq_addr   => count_order_inst_bus_wreq_addr,
      bus_wreq_len    => count_order_inst_bus_wreq_len,
      bus_wdat_valid  => count_order_inst_bus_wdat_valid,
      bus_wdat_ready  => count_order_inst_bus_wdat_ready,
      bus_wdat_data   => count_order_inst_bus_wdat_data,
      bus_wdat_strobe => count_order_inst_bus_wdat_strobe,
      bus_wdat_last   => count_order_inst_bus_wdat_last,
      in_valid        => count_order_inst_in_valid,
      in_ready        => count_order_inst_in_ready,
      in_data         => count_order_inst_in_data,
      in_dvalid       => count_order_inst_in_dvalid,
      in_last         => count_order_inst_in_last
    );

  l_returnflag_o_bus_wreq_valid      <= returnflag_o_inst_bus_wreq_valid;
  returnflag_o_inst_bus_wreq_ready   <= l_returnflag_o_bus_wreq_ready;
  l_returnflag_o_bus_wreq_addr       <= returnflag_o_inst_bus_wreq_addr;
  l_returnflag_o_bus_wreq_len        <= returnflag_o_inst_bus_wreq_len;
  l_returnflag_o_bus_wdat_valid      <= returnflag_o_inst_bus_wdat_valid;
  returnflag_o_inst_bus_wdat_ready   <= l_returnflag_o_bus_wdat_ready;
  l_returnflag_o_bus_wdat_data       <= returnflag_o_inst_bus_wdat_data;
  l_returnflag_o_bus_wdat_strobe     <= returnflag_o_inst_bus_wdat_strobe;
  l_returnflag_o_bus_wdat_last       <= returnflag_o_inst_bus_wdat_last;

  l_returnflag_o_unl_valid           <= returnflag_o_inst_unl_valid;
  returnflag_o_inst_unl_ready        <= l_returnflag_o_unl_ready;
  l_returnflag_o_unl_tag             <= returnflag_o_inst_unl_tag;

  l_linestatus_o_bus_wreq_valid      <= linestatus_o_inst_bus_wreq_valid;
  linestatus_o_inst_bus_wreq_ready   <= l_linestatus_o_bus_wreq_ready;
  l_linestatus_o_bus_wreq_addr       <= linestatus_o_inst_bus_wreq_addr;
  l_linestatus_o_bus_wreq_len        <= linestatus_o_inst_bus_wreq_len;
  l_linestatus_o_bus_wdat_valid      <= linestatus_o_inst_bus_wdat_valid;
  linestatus_o_inst_bus_wdat_ready   <= l_linestatus_o_bus_wdat_ready;
  l_linestatus_o_bus_wdat_data       <= linestatus_o_inst_bus_wdat_data;
  l_linestatus_o_bus_wdat_strobe     <= linestatus_o_inst_bus_wdat_strobe;
  l_linestatus_o_bus_wdat_last       <= linestatus_o_inst_bus_wdat_last;

  l_linestatus_o_unl_valid           <= linestatus_o_inst_unl_valid;
  linestatus_o_inst_unl_ready        <= l_linestatus_o_unl_ready;
  l_linestatus_o_unl_tag             <= linestatus_o_inst_unl_tag;

  l_sum_qty_bus_wreq_valid           <= sum_qty_inst_bus_wreq_valid;
  sum_qty_inst_bus_wreq_ready        <= l_sum_qty_bus_wreq_ready;
  l_sum_qty_bus_wreq_addr            <= sum_qty_inst_bus_wreq_addr;
  l_sum_qty_bus_wreq_len             <= sum_qty_inst_bus_wreq_len;
  l_sum_qty_bus_wdat_valid           <= sum_qty_inst_bus_wdat_valid;
  sum_qty_inst_bus_wdat_ready        <= l_sum_qty_bus_wdat_ready;
  l_sum_qty_bus_wdat_data            <= sum_qty_inst_bus_wdat_data;
  l_sum_qty_bus_wdat_strobe          <= sum_qty_inst_bus_wdat_strobe;
  l_sum_qty_bus_wdat_last            <= sum_qty_inst_bus_wdat_last;

  l_sum_qty_unl_valid                <= sum_qty_inst_unl_valid;
  sum_qty_inst_unl_ready             <= l_sum_qty_unl_ready;
  l_sum_qty_unl_tag                  <= sum_qty_inst_unl_tag;

  l_sum_base_price_bus_wreq_valid    <= sum_base_price_inst_bus_wreq_valid;
  sum_base_price_inst_bus_wreq_ready <= l_sum_base_price_bus_wreq_ready;
  l_sum_base_price_bus_wreq_addr     <= sum_base_price_inst_bus_wreq_addr;
  l_sum_base_price_bus_wreq_len      <= sum_base_price_inst_bus_wreq_len;
  l_sum_base_price_bus_wdat_valid    <= sum_base_price_inst_bus_wdat_valid;
  sum_base_price_inst_bus_wdat_ready <= l_sum_base_price_bus_wdat_ready;
  l_sum_base_price_bus_wdat_data     <= sum_base_price_inst_bus_wdat_data;
  l_sum_base_price_bus_wdat_strobe   <= sum_base_price_inst_bus_wdat_strobe;
  l_sum_base_price_bus_wdat_last     <= sum_base_price_inst_bus_wdat_last;

  l_sum_base_price_unl_valid         <= sum_base_price_inst_unl_valid;
  sum_base_price_inst_unl_ready      <= l_sum_base_price_unl_ready;
  l_sum_base_price_unl_tag           <= sum_base_price_inst_unl_tag;

  l_sum_disc_price_bus_wreq_valid    <= sum_disc_price_inst_bus_wreq_valid;
  sum_disc_price_inst_bus_wreq_ready <= l_sum_disc_price_bus_wreq_ready;
  l_sum_disc_price_bus_wreq_addr     <= sum_disc_price_inst_bus_wreq_addr;
  l_sum_disc_price_bus_wreq_len      <= sum_disc_price_inst_bus_wreq_len;
  l_sum_disc_price_bus_wdat_valid    <= sum_disc_price_inst_bus_wdat_valid;
  sum_disc_price_inst_bus_wdat_ready <= l_sum_disc_price_bus_wdat_ready;
  l_sum_disc_price_bus_wdat_data     <= sum_disc_price_inst_bus_wdat_data;
  l_sum_disc_price_bus_wdat_strobe   <= sum_disc_price_inst_bus_wdat_strobe;
  l_sum_disc_price_bus_wdat_last     <= sum_disc_price_inst_bus_wdat_last;

  l_sum_disc_price_unl_valid         <= sum_disc_price_inst_unl_valid;
  sum_disc_price_inst_unl_ready      <= l_sum_disc_price_unl_ready;
  l_sum_disc_price_unl_tag           <= sum_disc_price_inst_unl_tag;

  l_sum_charge_bus_wreq_valid        <= sum_charge_inst_bus_wreq_valid;
  sum_charge_inst_bus_wreq_ready     <= l_sum_charge_bus_wreq_ready;
  l_sum_charge_bus_wreq_addr         <= sum_charge_inst_bus_wreq_addr;
  l_sum_charge_bus_wreq_len          <= sum_charge_inst_bus_wreq_len;
  l_sum_charge_bus_wdat_valid        <= sum_charge_inst_bus_wdat_valid;
  sum_charge_inst_bus_wdat_ready     <= l_sum_charge_bus_wdat_ready;
  l_sum_charge_bus_wdat_data         <= sum_charge_inst_bus_wdat_data;
  l_sum_charge_bus_wdat_strobe       <= sum_charge_inst_bus_wdat_strobe;
  l_sum_charge_bus_wdat_last         <= sum_charge_inst_bus_wdat_last;

  l_sum_charge_unl_valid             <= sum_charge_inst_unl_valid;
  sum_charge_inst_unl_ready          <= l_sum_charge_unl_ready;
  l_sum_charge_unl_tag               <= sum_charge_inst_unl_tag;

  l_avg_qty_bus_wreq_valid           <= avg_qty_inst_bus_wreq_valid;
  avg_qty_inst_bus_wreq_ready        <= l_avg_qty_bus_wreq_ready;
  l_avg_qty_bus_wreq_addr            <= avg_qty_inst_bus_wreq_addr;
  l_avg_qty_bus_wreq_len             <= avg_qty_inst_bus_wreq_len;
  l_avg_qty_bus_wdat_valid           <= avg_qty_inst_bus_wdat_valid;
  avg_qty_inst_bus_wdat_ready        <= l_avg_qty_bus_wdat_ready;
  l_avg_qty_bus_wdat_data            <= avg_qty_inst_bus_wdat_data;
  l_avg_qty_bus_wdat_strobe          <= avg_qty_inst_bus_wdat_strobe;
  l_avg_qty_bus_wdat_last            <= avg_qty_inst_bus_wdat_last;

  l_avg_qty_unl_valid                <= avg_qty_inst_unl_valid;
  avg_qty_inst_unl_ready             <= l_avg_qty_unl_ready;
  l_avg_qty_unl_tag                  <= avg_qty_inst_unl_tag;

  l_avg_price_bus_wreq_valid         <= avg_price_inst_bus_wreq_valid;
  avg_price_inst_bus_wreq_ready      <= l_avg_price_bus_wreq_ready;
  l_avg_price_bus_wreq_addr          <= avg_price_inst_bus_wreq_addr;
  l_avg_price_bus_wreq_len           <= avg_price_inst_bus_wreq_len;
  l_avg_price_bus_wdat_valid         <= avg_price_inst_bus_wdat_valid;
  avg_price_inst_bus_wdat_ready      <= l_avg_price_bus_wdat_ready;
  l_avg_price_bus_wdat_data          <= avg_price_inst_bus_wdat_data;
  l_avg_price_bus_wdat_strobe        <= avg_price_inst_bus_wdat_strobe;
  l_avg_price_bus_wdat_last          <= avg_price_inst_bus_wdat_last;

  l_avg_price_unl_valid              <= avg_price_inst_unl_valid;
  avg_price_inst_unl_ready           <= l_avg_price_unl_ready;
  l_avg_price_unl_tag                <= avg_price_inst_unl_tag;

  l_avg_disc_bus_wreq_valid          <= avg_disc_inst_bus_wreq_valid;
  avg_disc_inst_bus_wreq_ready       <= l_avg_disc_bus_wreq_ready;
  l_avg_disc_bus_wreq_addr           <= avg_disc_inst_bus_wreq_addr;
  l_avg_disc_bus_wreq_len            <= avg_disc_inst_bus_wreq_len;
  l_avg_disc_bus_wdat_valid          <= avg_disc_inst_bus_wdat_valid;
  avg_disc_inst_bus_wdat_ready       <= l_avg_disc_bus_wdat_ready;
  l_avg_disc_bus_wdat_data           <= avg_disc_inst_bus_wdat_data;
  l_avg_disc_bus_wdat_strobe         <= avg_disc_inst_bus_wdat_strobe;
  l_avg_disc_bus_wdat_last           <= avg_disc_inst_bus_wdat_last;

  l_avg_disc_unl_valid               <= avg_disc_inst_unl_valid;
  avg_disc_inst_unl_ready            <= l_avg_disc_unl_ready;
  l_avg_disc_unl_tag                 <= avg_disc_inst_unl_tag;

  l_count_order_bus_wreq_valid       <= count_order_inst_bus_wreq_valid;
  count_order_inst_bus_wreq_ready    <= l_count_order_bus_wreq_ready;
  l_count_order_bus_wreq_addr        <= count_order_inst_bus_wreq_addr;
  l_count_order_bus_wreq_len         <= count_order_inst_bus_wreq_len;
  l_count_order_bus_wdat_valid       <= count_order_inst_bus_wdat_valid;
  count_order_inst_bus_wdat_ready    <= l_count_order_bus_wdat_ready;
  l_count_order_bus_wdat_data        <= count_order_inst_bus_wdat_data;
  l_count_order_bus_wdat_strobe      <= count_order_inst_bus_wdat_strobe;
  l_count_order_bus_wdat_last        <= count_order_inst_bus_wdat_last;

  l_count_order_unl_valid            <= count_order_inst_unl_valid;
  count_order_inst_unl_ready         <= l_count_order_unl_ready;
  l_count_order_unl_tag              <= count_order_inst_unl_tag;

  returnflag_o_inst_cmd_valid             <= l_returnflag_o_cmd_valid;
  l_returnflag_o_cmd_ready                <= returnflag_o_inst_cmd_ready;
  returnflag_o_inst_cmd_firstIdx          <= l_returnflag_o_cmd_firstIdx;
  returnflag_o_inst_cmd_lastIdx           <= l_returnflag_o_cmd_lastIdx;
  returnflag_o_inst_cmd_ctrl              <= l_returnflag_o_cmd_ctrl;
  returnflag_o_inst_cmd_tag               <= l_returnflag_o_cmd_tag;

  returnflag_o_inst_in_valid(0)           <= l_returnflag_o_valid;
  returnflag_o_inst_in_valid(1)           <= l_returnflag_o_chars_valid;
  l_returnflag_o_ready                    <= returnflag_o_inst_in_ready(0);
  l_returnflag_o_chars_ready              <= returnflag_o_inst_in_ready(1);
  returnflag_o_inst_in_data(31 downto 0)  <= l_returnflag_o_length;
  returnflag_o_inst_in_data(32 downto 32) <= l_returnflag_o_count;
  returnflag_o_inst_in_data(40 downto 33) <= l_returnflag_o_chars;
  returnflag_o_inst_in_data(41 downto 41) <= l_returnflag_o_chars_count;
  returnflag_o_inst_in_dvalid(0)          <= l_returnflag_o_dvalid;
  returnflag_o_inst_in_dvalid(1)          <= l_returnflag_o_chars_dvalid;
  returnflag_o_inst_in_last(0)            <= l_returnflag_o_last;
  returnflag_o_inst_in_last(1)            <= l_returnflag_o_chars_last;

  linestatus_o_inst_cmd_valid             <= l_linestatus_o_cmd_valid;
  l_linestatus_o_cmd_ready                <= linestatus_o_inst_cmd_ready;
  linestatus_o_inst_cmd_firstIdx          <= l_linestatus_o_cmd_firstIdx;
  linestatus_o_inst_cmd_lastIdx           <= l_linestatus_o_cmd_lastIdx;
  linestatus_o_inst_cmd_ctrl              <= l_linestatus_o_cmd_ctrl;
  linestatus_o_inst_cmd_tag               <= l_linestatus_o_cmd_tag;

  linestatus_o_inst_in_valid(0)           <= l_linestatus_o_valid;
  linestatus_o_inst_in_valid(1)           <= l_linestatus_o_chars_valid;
  l_linestatus_o_ready                    <= linestatus_o_inst_in_ready(0);
  l_linestatus_o_chars_ready              <= linestatus_o_inst_in_ready(1);
  linestatus_o_inst_in_data(31 downto 0)  <= l_linestatus_o_length;
  linestatus_o_inst_in_data(32 downto 32) <= l_linestatus_o_count;
  linestatus_o_inst_in_data(40 downto 33) <= l_linestatus_o_chars;
  linestatus_o_inst_in_data(41 downto 41) <= l_linestatus_o_chars_count;
  linestatus_o_inst_in_dvalid(0)          <= l_linestatus_o_dvalid;
  linestatus_o_inst_in_dvalid(1)          <= l_linestatus_o_chars_dvalid;
  linestatus_o_inst_in_last(0)            <= l_linestatus_o_last;
  linestatus_o_inst_in_last(1)            <= l_linestatus_o_chars_last;

  sum_qty_inst_cmd_valid                  <= l_sum_qty_cmd_valid;
  l_sum_qty_cmd_ready                     <= sum_qty_inst_cmd_ready;
  sum_qty_inst_cmd_firstIdx               <= l_sum_qty_cmd_firstIdx;
  sum_qty_inst_cmd_lastIdx                <= l_sum_qty_cmd_lastIdx;
  sum_qty_inst_cmd_ctrl                   <= l_sum_qty_cmd_ctrl;
  sum_qty_inst_cmd_tag                    <= l_sum_qty_cmd_tag;

  sum_qty_inst_in_valid(0)                <= l_sum_qty_valid;
  l_sum_qty_ready                         <= sum_qty_inst_in_ready(0);
  sum_qty_inst_in_data                    <= l_sum_qty;
  sum_qty_inst_in_dvalid(0)               <= l_sum_qty_dvalid;
  sum_qty_inst_in_last(0)                 <= l_sum_qty_last;

  sum_base_price_inst_cmd_valid           <= l_sum_base_price_cmd_valid;
  l_sum_base_price_cmd_ready              <= sum_base_price_inst_cmd_ready;
  sum_base_price_inst_cmd_firstIdx        <= l_sum_base_price_cmd_firstIdx;
  sum_base_price_inst_cmd_lastIdx         <= l_sum_base_price_cmd_lastIdx;
  sum_base_price_inst_cmd_ctrl            <= l_sum_base_price_cmd_ctrl;
  sum_base_price_inst_cmd_tag             <= l_sum_base_price_cmd_tag;

  sum_base_price_inst_in_valid(0)         <= l_sum_base_price_valid;
  l_sum_base_price_ready                  <= sum_base_price_inst_in_ready(0);
  sum_base_price_inst_in_data             <= l_sum_base_price;
  sum_base_price_inst_in_dvalid(0)        <= l_sum_base_price_dvalid;
  sum_base_price_inst_in_last(0)          <= l_sum_base_price_last;

  sum_disc_price_inst_cmd_valid           <= l_sum_disc_price_cmd_valid;
  l_sum_disc_price_cmd_ready              <= sum_disc_price_inst_cmd_ready;
  sum_disc_price_inst_cmd_firstIdx        <= l_sum_disc_price_cmd_firstIdx;
  sum_disc_price_inst_cmd_lastIdx         <= l_sum_disc_price_cmd_lastIdx;
  sum_disc_price_inst_cmd_ctrl            <= l_sum_disc_price_cmd_ctrl;
  sum_disc_price_inst_cmd_tag             <= l_sum_disc_price_cmd_tag;

  sum_disc_price_inst_in_valid(0)         <= l_sum_disc_price_valid;
  l_sum_disc_price_ready                  <= sum_disc_price_inst_in_ready(0);
  sum_disc_price_inst_in_data             <= l_sum_disc_price;
  sum_disc_price_inst_in_dvalid(0)        <= l_sum_disc_price_dvalid;
  sum_disc_price_inst_in_last(0)          <= l_sum_disc_price_last;

  sum_charge_inst_cmd_valid               <= l_sum_charge_cmd_valid;
  l_sum_charge_cmd_ready                  <= sum_charge_inst_cmd_ready;
  sum_charge_inst_cmd_firstIdx            <= l_sum_charge_cmd_firstIdx;
  sum_charge_inst_cmd_lastIdx             <= l_sum_charge_cmd_lastIdx;
  sum_charge_inst_cmd_ctrl                <= l_sum_charge_cmd_ctrl;
  sum_charge_inst_cmd_tag                 <= l_sum_charge_cmd_tag;

  sum_charge_inst_in_valid(0)             <= l_sum_charge_valid;
  l_sum_charge_ready                      <= sum_charge_inst_in_ready(0);
  sum_charge_inst_in_data                 <= l_sum_charge;
  sum_charge_inst_in_dvalid(0)            <= l_sum_charge_dvalid;
  sum_charge_inst_in_last(0)              <= l_sum_charge_last;

  avg_qty_inst_cmd_valid                  <= l_avg_qty_cmd_valid;
  l_avg_qty_cmd_ready                     <= avg_qty_inst_cmd_ready;
  avg_qty_inst_cmd_firstIdx               <= l_avg_qty_cmd_firstIdx;
  avg_qty_inst_cmd_lastIdx                <= l_avg_qty_cmd_lastIdx;
  avg_qty_inst_cmd_ctrl                   <= l_avg_qty_cmd_ctrl;
  avg_qty_inst_cmd_tag                    <= l_avg_qty_cmd_tag;

  avg_qty_inst_in_valid(0)                <= l_avg_qty_valid;
  l_avg_qty_ready                         <= avg_qty_inst_in_ready(0);
  avg_qty_inst_in_data                    <= l_avg_qty;
  avg_qty_inst_in_dvalid(0)               <= l_avg_qty_dvalid;
  avg_qty_inst_in_last(0)                 <= l_avg_qty_last;

  avg_price_inst_cmd_valid                <= l_avg_price_cmd_valid;
  l_avg_price_cmd_ready                   <= avg_price_inst_cmd_ready;
  avg_price_inst_cmd_firstIdx             <= l_avg_price_cmd_firstIdx;
  avg_price_inst_cmd_lastIdx              <= l_avg_price_cmd_lastIdx;
  avg_price_inst_cmd_ctrl                 <= l_avg_price_cmd_ctrl;
  avg_price_inst_cmd_tag                  <= l_avg_price_cmd_tag;

  avg_price_inst_in_valid(0)              <= l_avg_price_valid;
  l_avg_price_ready                       <= avg_price_inst_in_ready(0);
  avg_price_inst_in_data                  <= l_avg_price;
  avg_price_inst_in_dvalid(0)             <= l_avg_price_dvalid;
  avg_price_inst_in_last(0)               <= l_avg_price_last;

  avg_disc_inst_cmd_valid                 <= l_avg_disc_cmd_valid;
  l_avg_disc_cmd_ready                    <= avg_disc_inst_cmd_ready;
  avg_disc_inst_cmd_firstIdx              <= l_avg_disc_cmd_firstIdx;
  avg_disc_inst_cmd_lastIdx               <= l_avg_disc_cmd_lastIdx;
  avg_disc_inst_cmd_ctrl                  <= l_avg_disc_cmd_ctrl;
  avg_disc_inst_cmd_tag                   <= l_avg_disc_cmd_tag;

  avg_disc_inst_in_valid(0)               <= l_avg_disc_valid;
  l_avg_disc_ready                        <= avg_disc_inst_in_ready(0);
  avg_disc_inst_in_data                   <= l_avg_disc;
  avg_disc_inst_in_dvalid(0)              <= l_avg_disc_dvalid;
  avg_disc_inst_in_last(0)                <= l_avg_disc_last;

  count_order_inst_cmd_valid              <= l_count_order_cmd_valid;
  l_count_order_cmd_ready                 <= count_order_inst_cmd_ready;
  count_order_inst_cmd_firstIdx           <= l_count_order_cmd_firstIdx;
  count_order_inst_cmd_lastIdx            <= l_count_order_cmd_lastIdx;
  count_order_inst_cmd_ctrl               <= l_count_order_cmd_ctrl;
  count_order_inst_cmd_tag                <= l_count_order_cmd_tag;

  count_order_inst_in_valid(0)            <= l_count_order_valid;
  l_count_order_ready                     <= count_order_inst_in_ready(0);
  count_order_inst_in_data                <= l_count_order;
  count_order_inst_in_dvalid(0)           <= l_count_order_dvalid;
  count_order_inst_in_last(0)             <= l_count_order_last;

end architecture;
