-- Copyright 2018-2019 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
-- This file was generated by Fletchgen. Modify this file at your own risk.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.Array_pkg.all;

entity PriceSummary_l is
  generic (
    INDEX_WIDTH                         : integer := 32;
    TAG_WIDTH                           : integer := 1;
    L_QUANTITY_BUS_ADDR_WIDTH           : integer := 64;
    L_QUANTITY_BUS_DATA_WIDTH           : integer := 512;
    L_QUANTITY_BUS_LEN_WIDTH            : integer := 8;
    L_QUANTITY_BUS_BURST_STEP_LEN       : integer := 1;
    L_QUANTITY_BUS_BURST_MAX_LEN        : integer := 16;
    L_EXTENDEDPRICE_BUS_ADDR_WIDTH      : integer := 64;
    L_EXTENDEDPRICE_BUS_DATA_WIDTH      : integer := 512;
    L_EXTENDEDPRICE_BUS_LEN_WIDTH       : integer := 8;
    L_EXTENDEDPRICE_BUS_BURST_STEP_LEN  : integer := 1;
    L_EXTENDEDPRICE_BUS_BURST_MAX_LEN   : integer := 16;
    L_DISCOUNT_BUS_ADDR_WIDTH           : integer := 64;
    L_DISCOUNT_BUS_DATA_WIDTH           : integer := 512;
    L_DISCOUNT_BUS_LEN_WIDTH            : integer := 8;
    L_DISCOUNT_BUS_BURST_STEP_LEN       : integer := 1;
    L_DISCOUNT_BUS_BURST_MAX_LEN        : integer := 16;
    L_TAX_BUS_ADDR_WIDTH                : integer := 64;
    L_TAX_BUS_DATA_WIDTH                : integer := 512;
    L_TAX_BUS_LEN_WIDTH                 : integer := 8;
    L_TAX_BUS_BURST_STEP_LEN            : integer := 1;
    L_TAX_BUS_BURST_MAX_LEN             : integer := 16;
    L_RETURNFLAG_BUS_ADDR_WIDTH         : integer := 64;
    L_RETURNFLAG_BUS_DATA_WIDTH         : integer := 512;
    L_RETURNFLAG_BUS_LEN_WIDTH          : integer := 8;
    L_RETURNFLAG_BUS_BURST_STEP_LEN     : integer := 1;
    L_RETURNFLAG_BUS_BURST_MAX_LEN      : integer := 16;
    L_LINESTATUS_BUS_ADDR_WIDTH         : integer := 64;
    L_LINESTATUS_BUS_DATA_WIDTH         : integer := 512;
    L_LINESTATUS_BUS_LEN_WIDTH          : integer := 8;
    L_LINESTATUS_BUS_BURST_STEP_LEN     : integer := 1;
    L_LINESTATUS_BUS_BURST_MAX_LEN      : integer := 16;
    L_SHIPDATE_BUS_ADDR_WIDTH           : integer := 64;
    L_SHIPDATE_BUS_DATA_WIDTH           : integer := 512;
    L_SHIPDATE_BUS_LEN_WIDTH            : integer := 8;
    L_SHIPDATE_BUS_BURST_STEP_LEN       : integer := 1;
    L_SHIPDATE_BUS_BURST_MAX_LEN        : integer := 16;
    L_RETURNFLAG_O_BUS_ADDR_WIDTH       : integer := 64;
    L_RETURNFLAG_O_BUS_DATA_WIDTH       : integer := 512;
    L_RETURNFLAG_O_BUS_LEN_WIDTH        : integer := 8;
    L_RETURNFLAG_O_BUS_BURST_STEP_LEN   : integer := 1;
    L_RETURNFLAG_O_BUS_BURST_MAX_LEN    : integer := 16;
    L_LINESTATUS_O_BUS_ADDR_WIDTH       : integer := 64;
    L_LINESTATUS_O_BUS_DATA_WIDTH       : integer := 512;
    L_LINESTATUS_O_BUS_LEN_WIDTH        : integer := 8;
    L_LINESTATUS_O_BUS_BURST_STEP_LEN   : integer := 1;
    L_LINESTATUS_O_BUS_BURST_MAX_LEN    : integer := 16;
    L_SUM_QTY_BUS_ADDR_WIDTH            : integer := 64;
    L_SUM_QTY_BUS_DATA_WIDTH            : integer := 512;
    L_SUM_QTY_BUS_LEN_WIDTH             : integer := 8;
    L_SUM_QTY_BUS_BURST_STEP_LEN        : integer := 1;
    L_SUM_QTY_BUS_BURST_MAX_LEN         : integer := 16;
    L_SUM_BASE_PRICE_BUS_ADDR_WIDTH     : integer := 64;
    L_SUM_BASE_PRICE_BUS_DATA_WIDTH     : integer := 512;
    L_SUM_BASE_PRICE_BUS_LEN_WIDTH      : integer := 8;
    L_SUM_BASE_PRICE_BUS_BURST_STEP_LEN : integer := 1;
    L_SUM_BASE_PRICE_BUS_BURST_MAX_LEN  : integer := 16;
    L_SUM_DISC_PRICE_BUS_ADDR_WIDTH     : integer := 64;
    L_SUM_DISC_PRICE_BUS_DATA_WIDTH     : integer := 512;
    L_SUM_DISC_PRICE_BUS_LEN_WIDTH      : integer := 8;
    L_SUM_DISC_PRICE_BUS_BURST_STEP_LEN : integer := 1;
    L_SUM_DISC_PRICE_BUS_BURST_MAX_LEN  : integer := 16;
    L_SUM_CHARGE_BUS_ADDR_WIDTH         : integer := 64;
    L_SUM_CHARGE_BUS_DATA_WIDTH         : integer := 512;
    L_SUM_CHARGE_BUS_LEN_WIDTH          : integer := 8;
    L_SUM_CHARGE_BUS_BURST_STEP_LEN     : integer := 1;
    L_SUM_CHARGE_BUS_BURST_MAX_LEN      : integer := 16;
    L_AVG_QTY_BUS_ADDR_WIDTH            : integer := 64;
    L_AVG_QTY_BUS_DATA_WIDTH            : integer := 512;
    L_AVG_QTY_BUS_LEN_WIDTH             : integer := 8;
    L_AVG_QTY_BUS_BURST_STEP_LEN        : integer := 1;
    L_AVG_QTY_BUS_BURST_MAX_LEN         : integer := 16;
    L_AVG_PRICE_BUS_ADDR_WIDTH          : integer := 64;
    L_AVG_PRICE_BUS_DATA_WIDTH          : integer := 512;
    L_AVG_PRICE_BUS_LEN_WIDTH           : integer := 8;
    L_AVG_PRICE_BUS_BURST_STEP_LEN      : integer := 1;
    L_AVG_PRICE_BUS_BURST_MAX_LEN       : integer := 16;
    L_AVG_DISC_BUS_ADDR_WIDTH           : integer := 64;
    L_AVG_DISC_BUS_DATA_WIDTH           : integer := 512;
    L_AVG_DISC_BUS_LEN_WIDTH            : integer := 8;
    L_AVG_DISC_BUS_BURST_STEP_LEN       : integer := 1;
    L_AVG_DISC_BUS_BURST_MAX_LEN        : integer := 16;
    L_COUNT_ORDER_BUS_ADDR_WIDTH        : integer := 64;
    L_COUNT_ORDER_BUS_DATA_WIDTH        : integer := 512;
    L_COUNT_ORDER_BUS_LEN_WIDTH         : integer := 8;
    L_COUNT_ORDER_BUS_BURST_STEP_LEN    : integer := 1;
    L_COUNT_ORDER_BUS_BURST_MAX_LEN     : integer := 16
  );
  port (
    bcd_clk                          : in std_logic;
    bcd_reset                        : in std_logic;
    kcd_clk                          : in std_logic;
    kcd_reset                        : in std_logic;
    l_quantity_valid                 : out std_logic;
    l_quantity_ready                 : in std_logic;
    l_quantity_dvalid                : out std_logic;
    l_quantity_last                  : out std_logic;
    l_quantity                       : out std_logic_vector(63 downto 0);
    l_quantity_bus_rreq_valid        : out std_logic;
    l_quantity_bus_rreq_ready        : in std_logic;
    l_quantity_bus_rreq_addr         : out std_logic_vector(L_QUANTITY_BUS_ADDR_WIDTH - 1 downto 0);
    l_quantity_bus_rreq_len          : out std_logic_vector(L_QUANTITY_BUS_LEN_WIDTH - 1 downto 0);
    l_quantity_bus_rdat_valid        : in std_logic;
    l_quantity_bus_rdat_ready        : out std_logic;
    l_quantity_bus_rdat_data         : in std_logic_vector(L_QUANTITY_BUS_DATA_WIDTH - 1 downto 0);
    l_quantity_bus_rdat_last         : in std_logic;
    l_quantity_cmd_valid             : in std_logic;
    l_quantity_cmd_ready             : out std_logic;
    l_quantity_cmd_firstIdx          : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    l_quantity_cmd_lastIdx           : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    l_quantity_cmd_ctrl              : in std_logic_vector(L_QUANTITY_BUS_ADDR_WIDTH - 1 downto 0);
    l_quantity_cmd_tag               : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    l_quantity_unl_valid             : out std_logic;
    l_quantity_unl_ready             : in std_logic;
    l_quantity_unl_tag               : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    l_extendedprice_valid            : out std_logic;
    l_extendedprice_ready            : in std_logic;
    l_extendedprice_dvalid           : out std_logic;
    l_extendedprice_last             : out std_logic;
    l_extendedprice                  : out std_logic_vector(63 downto 0);
    l_extendedprice_bus_rreq_valid   : out std_logic;
    l_extendedprice_bus_rreq_ready   : in std_logic;
    l_extendedprice_bus_rreq_addr    : out std_logic_vector(L_EXTENDEDPRICE_BUS_ADDR_WIDTH - 1 downto 0);
    l_extendedprice_bus_rreq_len     : out std_logic_vector(L_EXTENDEDPRICE_BUS_LEN_WIDTH - 1 downto 0);
    l_extendedprice_bus_rdat_valid   : in std_logic;
    l_extendedprice_bus_rdat_ready   : out std_logic;
    l_extendedprice_bus_rdat_data    : in std_logic_vector(L_EXTENDEDPRICE_BUS_DATA_WIDTH - 1 downto 0);
    l_extendedprice_bus_rdat_last    : in std_logic;
    l_extendedprice_cmd_valid        : in std_logic;
    l_extendedprice_cmd_ready        : out std_logic;
    l_extendedprice_cmd_firstIdx     : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    l_extendedprice_cmd_lastIdx      : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    l_extendedprice_cmd_ctrl         : in std_logic_vector(L_EXTENDEDPRICE_BUS_ADDR_WIDTH - 1 downto 0);
    l_extendedprice_cmd_tag          : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    l_extendedprice_unl_valid        : out std_logic;
    l_extendedprice_unl_ready        : in std_logic;
    l_extendedprice_unl_tag          : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    l_discount_valid                 : out std_logic;
    l_discount_ready                 : in std_logic;
    l_discount_dvalid                : out std_logic;
    l_discount_last                  : out std_logic;
    l_discount                       : out std_logic_vector(63 downto 0);
    l_discount_bus_rreq_valid        : out std_logic;
    l_discount_bus_rreq_ready        : in std_logic;
    l_discount_bus_rreq_addr         : out std_logic_vector(L_DISCOUNT_BUS_ADDR_WIDTH - 1 downto 0);
    l_discount_bus_rreq_len          : out std_logic_vector(L_DISCOUNT_BUS_LEN_WIDTH - 1 downto 0);
    l_discount_bus_rdat_valid        : in std_logic;
    l_discount_bus_rdat_ready        : out std_logic;
    l_discount_bus_rdat_data         : in std_logic_vector(L_DISCOUNT_BUS_DATA_WIDTH - 1 downto 0);
    l_discount_bus_rdat_last         : in std_logic;
    l_discount_cmd_valid             : in std_logic;
    l_discount_cmd_ready             : out std_logic;
    l_discount_cmd_firstIdx          : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    l_discount_cmd_lastIdx           : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    l_discount_cmd_ctrl              : in std_logic_vector(L_DISCOUNT_BUS_ADDR_WIDTH - 1 downto 0);
    l_discount_cmd_tag               : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    l_discount_unl_valid             : out std_logic;
    l_discount_unl_ready             : in std_logic;
    l_discount_unl_tag               : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    l_tax_valid                      : out std_logic;
    l_tax_ready                      : in std_logic;
    l_tax_dvalid                     : out std_logic;
    l_tax_last                       : out std_logic;
    l_tax                            : out std_logic_vector(63 downto 0);
    l_tax_bus_rreq_valid             : out std_logic;
    l_tax_bus_rreq_ready             : in std_logic;
    l_tax_bus_rreq_addr              : out std_logic_vector(L_TAX_BUS_ADDR_WIDTH - 1 downto 0);
    l_tax_bus_rreq_len               : out std_logic_vector(L_TAX_BUS_LEN_WIDTH - 1 downto 0);
    l_tax_bus_rdat_valid             : in std_logic;
    l_tax_bus_rdat_ready             : out std_logic;
    l_tax_bus_rdat_data              : in std_logic_vector(L_TAX_BUS_DATA_WIDTH - 1 downto 0);
    l_tax_bus_rdat_last              : in std_logic;
    l_tax_cmd_valid                  : in std_logic;
    l_tax_cmd_ready                  : out std_logic;
    l_tax_cmd_firstIdx               : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    l_tax_cmd_lastIdx                : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    l_tax_cmd_ctrl                   : in std_logic_vector(L_TAX_BUS_ADDR_WIDTH - 1 downto 0);
    l_tax_cmd_tag                    : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    l_tax_unl_valid                  : out std_logic;
    l_tax_unl_ready                  : in std_logic;
    l_tax_unl_tag                    : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    l_returnflag_valid               : out std_logic;
    l_returnflag_ready               : in std_logic;
    l_returnflag_dvalid              : out std_logic;
    l_returnflag_last                : out std_logic;
    l_returnflag_length              : out std_logic_vector(31 downto 0);
    l_returnflag_count               : out std_logic_vector(0 downto 0);
    l_returnflag_chars_valid         : out std_logic;
    l_returnflag_chars_ready         : in std_logic;
    l_returnflag_chars_dvalid        : out std_logic;
    l_returnflag_chars_last          : out std_logic;
    l_returnflag_chars               : out std_logic_vector(7 downto 0);
    l_returnflag_chars_count         : out std_logic_vector(0 downto 0);
    l_returnflag_bus_rreq_valid      : out std_logic;
    l_returnflag_bus_rreq_ready      : in std_logic;
    l_returnflag_bus_rreq_addr       : out std_logic_vector(L_RETURNFLAG_BUS_ADDR_WIDTH - 1 downto 0);
    l_returnflag_bus_rreq_len        : out std_logic_vector(L_RETURNFLAG_BUS_LEN_WIDTH - 1 downto 0);
    l_returnflag_bus_rdat_valid      : in std_logic;
    l_returnflag_bus_rdat_ready      : out std_logic;
    l_returnflag_bus_rdat_data       : in std_logic_vector(L_RETURNFLAG_BUS_DATA_WIDTH - 1 downto 0);
    l_returnflag_bus_rdat_last       : in std_logic;
    l_returnflag_cmd_valid           : in std_logic;
    l_returnflag_cmd_ready           : out std_logic;
    l_returnflag_cmd_firstIdx        : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    l_returnflag_cmd_lastIdx         : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    l_returnflag_cmd_ctrl            : in std_logic_vector(L_RETURNFLAG_BUS_ADDR_WIDTH * 2 - 1 downto 0);
    l_returnflag_cmd_tag             : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    l_returnflag_unl_valid           : out std_logic;
    l_returnflag_unl_ready           : in std_logic;
    l_returnflag_unl_tag             : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    l_linestatus_valid               : out std_logic;
    l_linestatus_ready               : in std_logic;
    l_linestatus_dvalid              : out std_logic;
    l_linestatus_last                : out std_logic;
    l_linestatus_length              : out std_logic_vector(31 downto 0);
    l_linestatus_count               : out std_logic_vector(0 downto 0);
    l_linestatus_chars_valid         : out std_logic;
    l_linestatus_chars_ready         : in std_logic;
    l_linestatus_chars_dvalid        : out std_logic;
    l_linestatus_chars_last          : out std_logic;
    l_linestatus_chars               : out std_logic_vector(7 downto 0);
    l_linestatus_chars_count         : out std_logic_vector(0 downto 0);
    l_linestatus_bus_rreq_valid      : out std_logic;
    l_linestatus_bus_rreq_ready      : in std_logic;
    l_linestatus_bus_rreq_addr       : out std_logic_vector(L_LINESTATUS_BUS_ADDR_WIDTH - 1 downto 0);
    l_linestatus_bus_rreq_len        : out std_logic_vector(L_LINESTATUS_BUS_LEN_WIDTH - 1 downto 0);
    l_linestatus_bus_rdat_valid      : in std_logic;
    l_linestatus_bus_rdat_ready      : out std_logic;
    l_linestatus_bus_rdat_data       : in std_logic_vector(L_LINESTATUS_BUS_DATA_WIDTH - 1 downto 0);
    l_linestatus_bus_rdat_last       : in std_logic;
    l_linestatus_cmd_valid           : in std_logic;
    l_linestatus_cmd_ready           : out std_logic;
    l_linestatus_cmd_firstIdx        : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    l_linestatus_cmd_lastIdx         : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    l_linestatus_cmd_ctrl            : in std_logic_vector(L_LINESTATUS_BUS_ADDR_WIDTH * 2 - 1 downto 0);
    l_linestatus_cmd_tag             : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    l_linestatus_unl_valid           : out std_logic;
    l_linestatus_unl_ready           : in std_logic;
    l_linestatus_unl_tag             : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    l_shipdate_valid                 : out std_logic;
    l_shipdate_ready                 : in std_logic;
    l_shipdate_dvalid                : out std_logic;
    l_shipdate_last                  : out std_logic;
    l_shipdate                       : out std_logic_vector(31 downto 0);
    l_shipdate_bus_rreq_valid        : out std_logic;
    l_shipdate_bus_rreq_ready        : in std_logic;
    l_shipdate_bus_rreq_addr         : out std_logic_vector(L_SHIPDATE_BUS_ADDR_WIDTH - 1 downto 0);
    l_shipdate_bus_rreq_len          : out std_logic_vector(L_SHIPDATE_BUS_LEN_WIDTH - 1 downto 0);
    l_shipdate_bus_rdat_valid        : in std_logic;
    l_shipdate_bus_rdat_ready        : out std_logic;
    l_shipdate_bus_rdat_data         : in std_logic_vector(L_SHIPDATE_BUS_DATA_WIDTH - 1 downto 0);
    l_shipdate_bus_rdat_last         : in std_logic;
    l_shipdate_cmd_valid             : in std_logic;
    l_shipdate_cmd_ready             : out std_logic;
    l_shipdate_cmd_firstIdx          : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    l_shipdate_cmd_lastIdx           : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    l_shipdate_cmd_ctrl              : in std_logic_vector(L_SHIPDATE_BUS_ADDR_WIDTH - 1 downto 0);
    l_shipdate_cmd_tag               : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    l_shipdate_unl_valid             : out std_logic;
    l_shipdate_unl_ready             : in std_logic;
    l_shipdate_unl_tag               : out std_logic_vector(TAG_WIDTH - 1 downto 0);

    l_returnflag_o_valid             : in std_logic;
    l_returnflag_o_ready             : out std_logic;
    l_returnflag_o_dvalid            : in std_logic;
    l_returnflag_o_last              : in std_logic;
    l_returnflag_o_length            : in std_logic_vector(31 downto 0);
    l_returnflag_o_count             : in std_logic_vector(0 downto 0);
    l_returnflag_o_chars_valid       : in std_logic;
    l_returnflag_o_chars_ready       : out std_logic;
    l_returnflag_o_chars_dvalid      : in std_logic;
    l_returnflag_o_chars_last        : in std_logic;
    l_returnflag_o_chars             : in std_logic_vector(7 downto 0);
    l_returnflag_o_chars_count       : in std_logic_vector(0 downto 0);
    l_returnflag_o_bus_wreq_valid    : out std_logic;
    l_returnflag_o_bus_wreq_ready    : in std_logic;
    l_returnflag_o_bus_wreq_addr     : out std_logic_vector(L_RETURNFLAG_O_BUS_ADDR_WIDTH - 1 downto 0);
    l_returnflag_o_bus_wreq_len      : out std_logic_vector(L_RETURNFLAG_O_BUS_LEN_WIDTH - 1 downto 0);
    l_returnflag_o_bus_wreq_last     : out std_logic;
    l_returnflag_o_bus_wdat_valid    : out std_logic;
    l_returnflag_o_bus_wdat_ready    : in std_logic;
    l_returnflag_o_bus_wdat_data     : out std_logic_vector(L_RETURNFLAG_O_BUS_DATA_WIDTH - 1 downto 0);
    l_returnflag_o_bus_wdat_strobe   : out std_logic_vector(L_RETURNFLAG_O_BUS_DATA_WIDTH/8 - 1 downto 0);
    l_returnflag_o_bus_wdat_last     : out std_logic;
    l_returnflag_o_bus_wrep_valid    : in std_logic;
    l_returnflag_o_bus_wrep_ready    : out std_logic;
    l_returnflag_o_bus_wrep_ok       : in std_logic;
    l_returnflag_o_cmd_valid         : in std_logic;
    l_returnflag_o_cmd_ready         : out std_logic;
    l_returnflag_o_cmd_firstIdx      : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    l_returnflag_o_cmd_lastIdx       : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    l_returnflag_o_cmd_ctrl          : in std_logic_vector(L_RETURNFLAG_O_BUS_ADDR_WIDTH * 2 - 1 downto 0);
    l_returnflag_o_cmd_tag           : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    l_returnflag_o_unl_valid         : out std_logic;
    l_returnflag_o_unl_ready         : in std_logic;
    l_returnflag_o_unl_tag           : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    l_linestatus_o_valid             : in std_logic;
    l_linestatus_o_ready             : out std_logic;
    l_linestatus_o_dvalid            : in std_logic;
    l_linestatus_o_last              : in std_logic;
    l_linestatus_o_length            : in std_logic_vector(31 downto 0);
    l_linestatus_o_count             : in std_logic_vector(0 downto 0);
    l_linestatus_o_chars_valid       : in std_logic;
    l_linestatus_o_chars_ready       : out std_logic;
    l_linestatus_o_chars_dvalid      : in std_logic;
    l_linestatus_o_chars_last        : in std_logic;
    l_linestatus_o_chars             : in std_logic_vector(7 downto 0);
    l_linestatus_o_chars_count       : in std_logic_vector(0 downto 0);
    l_linestatus_o_bus_wreq_valid    : out std_logic;
    l_linestatus_o_bus_wreq_ready    : in std_logic;
    l_linestatus_o_bus_wreq_addr     : out std_logic_vector(L_LINESTATUS_O_BUS_ADDR_WIDTH - 1 downto 0);
    l_linestatus_o_bus_wreq_len      : out std_logic_vector(L_LINESTATUS_O_BUS_LEN_WIDTH - 1 downto 0);
    l_linestatus_o_bus_wreq_last     : out std_logic;
    l_linestatus_o_bus_wdat_valid    : out std_logic;
    l_linestatus_o_bus_wdat_ready    : in std_logic;
    l_linestatus_o_bus_wdat_data     : out std_logic_vector(L_LINESTATUS_O_BUS_DATA_WIDTH - 1 downto 0);
    l_linestatus_o_bus_wdat_strobe   : out std_logic_vector(L_LINESTATUS_O_BUS_DATA_WIDTH/8 - 1 downto 0);
    l_linestatus_o_bus_wdat_last     : out std_logic;
    l_linestatus_o_bus_wrep_valid    : in std_logic;
    l_linestatus_o_bus_wrep_ready    : out std_logic;
    l_linestatus_o_bus_wrep_ok       : in std_logic;
    l_linestatus_o_cmd_valid         : in std_logic;
    l_linestatus_o_cmd_ready         : out std_logic;
    l_linestatus_o_cmd_firstIdx      : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    l_linestatus_o_cmd_lastIdx       : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    l_linestatus_o_cmd_ctrl          : in std_logic_vector(L_LINESTATUS_O_BUS_ADDR_WIDTH * 2 - 1 downto 0);
    l_linestatus_o_cmd_tag           : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    l_linestatus_o_unl_valid         : out std_logic;
    l_linestatus_o_unl_ready         : in std_logic;
    l_linestatus_o_unl_tag           : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    l_sum_qty_valid                  : in std_logic;
    l_sum_qty_ready                  : out std_logic;
    l_sum_qty_dvalid                 : in std_logic;
    l_sum_qty_last                   : in std_logic;
    l_sum_qty                        : in std_logic_vector(63 downto 0);
    l_sum_qty_bus_wreq_valid         : out std_logic;
    l_sum_qty_bus_wreq_ready         : in std_logic;
    l_sum_qty_bus_wreq_addr          : out std_logic_vector(L_SUM_QTY_BUS_ADDR_WIDTH - 1 downto 0);
    l_sum_qty_bus_wreq_len           : out std_logic_vector(L_SUM_QTY_BUS_LEN_WIDTH - 1 downto 0);
    l_sum_qty_bus_wreq_last          : out std_logic;
    l_sum_qty_bus_wdat_valid         : out std_logic;
    l_sum_qty_bus_wdat_ready         : in std_logic;
    l_sum_qty_bus_wdat_data          : out std_logic_vector(L_SUM_QTY_BUS_DATA_WIDTH - 1 downto 0);
    l_sum_qty_bus_wdat_strobe        : out std_logic_vector(L_SUM_QTY_BUS_DATA_WIDTH/8 - 1 downto 0);
    l_sum_qty_bus_wdat_last          : out std_logic;
    l_sum_qty_bus_wrep_valid         : in std_logic;
    l_sum_qty_bus_wrep_ready         : out std_logic;
    l_sum_qty_bus_wrep_ok            : in std_logic;
    l_sum_qty_cmd_valid              : in std_logic;
    l_sum_qty_cmd_ready              : out std_logic;
    l_sum_qty_cmd_firstIdx           : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    l_sum_qty_cmd_lastIdx            : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    l_sum_qty_cmd_ctrl               : in std_logic_vector(L_SUM_QTY_BUS_ADDR_WIDTH - 1 downto 0);
    l_sum_qty_cmd_tag                : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    l_sum_qty_unl_valid              : out std_logic;
    l_sum_qty_unl_ready              : in std_logic;
    l_sum_qty_unl_tag                : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    l_sum_base_price_valid           : in std_logic;
    l_sum_base_price_ready           : out std_logic;
    l_sum_base_price_dvalid          : in std_logic;
    l_sum_base_price_last            : in std_logic;
    l_sum_base_price                 : in std_logic_vector(63 downto 0);
    l_sum_base_price_bus_wreq_valid  : out std_logic;
    l_sum_base_price_bus_wreq_ready  : in std_logic;
    l_sum_base_price_bus_wreq_addr   : out std_logic_vector(L_SUM_BASE_PRICE_BUS_ADDR_WIDTH - 1 downto 0);
    l_sum_base_price_bus_wreq_len    : out std_logic_vector(L_SUM_BASE_PRICE_BUS_LEN_WIDTH - 1 downto 0);
    l_sum_base_price_bus_wreq_last   : out std_logic;
    l_sum_base_price_bus_wdat_valid  : out std_logic;
    l_sum_base_price_bus_wdat_ready  : in std_logic;
    l_sum_base_price_bus_wdat_data   : out std_logic_vector(L_SUM_BASE_PRICE_BUS_DATA_WIDTH - 1 downto 0);
    l_sum_base_price_bus_wdat_strobe : out std_logic_vector(L_SUM_BASE_PRICE_BUS_DATA_WIDTH/8 - 1 downto 0);
    l_sum_base_price_bus_wdat_last   : out std_logic;
    l_sum_base_price_bus_wrep_valid  : in std_logic;
    l_sum_base_price_bus_wrep_ready  : out std_logic;
    l_sum_base_price_bus_wrep_ok     : in std_logic;
    l_sum_base_price_cmd_valid       : in std_logic;
    l_sum_base_price_cmd_ready       : out std_logic;
    l_sum_base_price_cmd_firstIdx    : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    l_sum_base_price_cmd_lastIdx     : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    l_sum_base_price_cmd_ctrl        : in std_logic_vector(L_SUM_BASE_PRICE_BUS_ADDR_WIDTH - 1 downto 0);
    l_sum_base_price_cmd_tag         : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    l_sum_base_price_unl_valid       : out std_logic;
    l_sum_base_price_unl_ready       : in std_logic;
    l_sum_base_price_unl_tag         : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    l_sum_disc_price_valid           : in std_logic;
    l_sum_disc_price_ready           : out std_logic;
    l_sum_disc_price_dvalid          : in std_logic;
    l_sum_disc_price_last            : in std_logic;
    l_sum_disc_price                 : in std_logic_vector(63 downto 0);
    l_sum_disc_price_bus_wreq_valid  : out std_logic;
    l_sum_disc_price_bus_wreq_ready  : in std_logic;
    l_sum_disc_price_bus_wreq_addr   : out std_logic_vector(L_SUM_DISC_PRICE_BUS_ADDR_WIDTH - 1 downto 0);
    l_sum_disc_price_bus_wreq_len    : out std_logic_vector(L_SUM_DISC_PRICE_BUS_LEN_WIDTH - 1 downto 0);
    l_sum_disc_price_bus_wreq_last   : out std_logic;
    l_sum_disc_price_bus_wdat_valid  : out std_logic;
    l_sum_disc_price_bus_wdat_ready  : in std_logic;
    l_sum_disc_price_bus_wdat_data   : out std_logic_vector(L_SUM_DISC_PRICE_BUS_DATA_WIDTH - 1 downto 0);
    l_sum_disc_price_bus_wdat_strobe : out std_logic_vector(L_SUM_DISC_PRICE_BUS_DATA_WIDTH/8 - 1 downto 0);
    l_sum_disc_price_bus_wdat_last   : out std_logic;
    l_sum_disc_price_bus_wrep_valid  : in std_logic;
    l_sum_disc_price_bus_wrep_ready  : out std_logic;
    l_sum_disc_price_bus_wrep_ok     : in std_logic;
    l_sum_disc_price_cmd_valid       : in std_logic;
    l_sum_disc_price_cmd_ready       : out std_logic;
    l_sum_disc_price_cmd_firstIdx    : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    l_sum_disc_price_cmd_lastIdx     : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    l_sum_disc_price_cmd_ctrl        : in std_logic_vector(L_SUM_DISC_PRICE_BUS_ADDR_WIDTH - 1 downto 0);
    l_sum_disc_price_cmd_tag         : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    l_sum_disc_price_unl_valid       : out std_logic;
    l_sum_disc_price_unl_ready       : in std_logic;
    l_sum_disc_price_unl_tag         : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    l_sum_charge_valid               : in std_logic;
    l_sum_charge_ready               : out std_logic;
    l_sum_charge_dvalid              : in std_logic;
    l_sum_charge_last                : in std_logic;
    l_sum_charge                     : in std_logic_vector(63 downto 0);
    l_sum_charge_bus_wreq_valid      : out std_logic;
    l_sum_charge_bus_wreq_ready      : in std_logic;
    l_sum_charge_bus_wreq_addr       : out std_logic_vector(L_SUM_CHARGE_BUS_ADDR_WIDTH - 1 downto 0);
    l_sum_charge_bus_wreq_len        : out std_logic_vector(L_SUM_CHARGE_BUS_LEN_WIDTH - 1 downto 0);
    l_sum_charge_bus_wreq_last       : out std_logic;
    l_sum_charge_bus_wdat_valid      : out std_logic;
    l_sum_charge_bus_wdat_ready      : in std_logic;
    l_sum_charge_bus_wdat_data       : out std_logic_vector(L_SUM_CHARGE_BUS_DATA_WIDTH - 1 downto 0);
    l_sum_charge_bus_wdat_strobe     : out std_logic_vector(L_SUM_CHARGE_BUS_DATA_WIDTH/8 - 1 downto 0);
    l_sum_charge_bus_wdat_last       : out std_logic;
    l_sum_charge_bus_wrep_valid      : in std_logic;
    l_sum_charge_bus_wrep_ready      : out std_logic;
    l_sum_charge_bus_wrep_ok         : in std_logic;
    l_sum_charge_cmd_valid           : in std_logic;
    l_sum_charge_cmd_ready           : out std_logic;
    l_sum_charge_cmd_firstIdx        : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    l_sum_charge_cmd_lastIdx         : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    l_sum_charge_cmd_ctrl            : in std_logic_vector(L_SUM_CHARGE_BUS_ADDR_WIDTH - 1 downto 0);
    l_sum_charge_cmd_tag             : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    l_sum_charge_unl_valid           : out std_logic;
    l_sum_charge_unl_ready           : in std_logic;
    l_sum_charge_unl_tag             : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    l_avg_qty_valid                  : in std_logic;
    l_avg_qty_ready                  : out std_logic;
    l_avg_qty_dvalid                 : in std_logic;
    l_avg_qty_last                   : in std_logic;
    l_avg_qty                        : in std_logic_vector(63 downto 0);
    l_avg_qty_bus_wreq_valid         : out std_logic;
    l_avg_qty_bus_wreq_ready         : in std_logic;
    l_avg_qty_bus_wreq_addr          : out std_logic_vector(L_AVG_QTY_BUS_ADDR_WIDTH - 1 downto 0);
    l_avg_qty_bus_wreq_len           : out std_logic_vector(L_AVG_QTY_BUS_LEN_WIDTH - 1 downto 0);
    l_avg_qty_bus_wreq_last          : out std_logic;
    l_avg_qty_bus_wdat_valid         : out std_logic;
    l_avg_qty_bus_wdat_ready         : in std_logic;
    l_avg_qty_bus_wdat_data          : out std_logic_vector(L_AVG_QTY_BUS_DATA_WIDTH - 1 downto 0);
    l_avg_qty_bus_wdat_strobe        : out std_logic_vector(L_AVG_QTY_BUS_DATA_WIDTH/8 - 1 downto 0);
    l_avg_qty_bus_wdat_last          : out std_logic;
    l_avg_qty_bus_wrep_valid         : in std_logic;
    l_avg_qty_bus_wrep_ready         : out std_logic;
    l_avg_qty_bus_wrep_ok            : in std_logic;
    l_avg_qty_cmd_valid              : in std_logic;
    l_avg_qty_cmd_ready              : out std_logic;
    l_avg_qty_cmd_firstIdx           : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    l_avg_qty_cmd_lastIdx            : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    l_avg_qty_cmd_ctrl               : in std_logic_vector(L_AVG_QTY_BUS_ADDR_WIDTH - 1 downto 0);
    l_avg_qty_cmd_tag                : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    l_avg_qty_unl_valid              : out std_logic;
    l_avg_qty_unl_ready              : in std_logic;
    l_avg_qty_unl_tag                : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    l_avg_price_valid                : in std_logic;
    l_avg_price_ready                : out std_logic;
    l_avg_price_dvalid               : in std_logic;
    l_avg_price_last                 : in std_logic;
    l_avg_price                      : in std_logic_vector(63 downto 0);
    l_avg_price_bus_wreq_valid       : out std_logic;
    l_avg_price_bus_wreq_ready       : in std_logic;
    l_avg_price_bus_wreq_addr        : out std_logic_vector(L_AVG_PRICE_BUS_ADDR_WIDTH - 1 downto 0);
    l_avg_price_bus_wreq_len         : out std_logic_vector(L_AVG_PRICE_BUS_LEN_WIDTH - 1 downto 0);
    l_avg_price_bus_wreq_last        : out std_logic;
    l_avg_price_bus_wdat_valid       : out std_logic;
    l_avg_price_bus_wdat_ready       : in std_logic;
    l_avg_price_bus_wdat_data        : out std_logic_vector(L_AVG_PRICE_BUS_DATA_WIDTH - 1 downto 0);
    l_avg_price_bus_wdat_strobe      : out std_logic_vector(L_AVG_PRICE_BUS_DATA_WIDTH/8 - 1 downto 0);
    l_avg_price_bus_wdat_last        : out std_logic;
    l_avg_price_bus_wrep_valid       : in std_logic;
    l_avg_price_bus_wrep_ready       : out std_logic;
    l_avg_price_bus_wrep_ok          : in std_logic;
    l_avg_price_cmd_valid            : in std_logic;
    l_avg_price_cmd_ready            : out std_logic;
    l_avg_price_cmd_firstIdx         : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    l_avg_price_cmd_lastIdx          : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    l_avg_price_cmd_ctrl             : in std_logic_vector(L_AVG_PRICE_BUS_ADDR_WIDTH - 1 downto 0);
    l_avg_price_cmd_tag              : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    l_avg_price_unl_valid            : out std_logic;
    l_avg_price_unl_ready            : in std_logic;
    l_avg_price_unl_tag              : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    l_avg_disc_valid                 : in std_logic;
    l_avg_disc_ready                 : out std_logic;
    l_avg_disc_dvalid                : in std_logic;
    l_avg_disc_last                  : in std_logic;
    l_avg_disc                       : in std_logic_vector(63 downto 0);
    l_avg_disc_bus_wreq_valid        : out std_logic;
    l_avg_disc_bus_wreq_ready        : in std_logic;
    l_avg_disc_bus_wreq_addr         : out std_logic_vector(L_AVG_DISC_BUS_ADDR_WIDTH - 1 downto 0);
    l_avg_disc_bus_wreq_len          : out std_logic_vector(L_AVG_DISC_BUS_LEN_WIDTH - 1 downto 0);
    l_avg_disc_bus_wreq_last         : out std_logic;
    l_avg_disc_bus_wdat_valid        : out std_logic;
    l_avg_disc_bus_wdat_ready        : in std_logic;
    l_avg_disc_bus_wdat_data         : out std_logic_vector(L_AVG_DISC_BUS_DATA_WIDTH - 1 downto 0);
    l_avg_disc_bus_wdat_strobe       : out std_logic_vector(L_AVG_DISC_BUS_DATA_WIDTH/8 - 1 downto 0);
    l_avg_disc_bus_wdat_last         : out std_logic;
    l_avg_disc_bus_wrep_valid        : in std_logic;
    l_avg_disc_bus_wrep_ready        : out std_logic;
    l_avg_disc_bus_wrep_ok           : in std_logic;
    l_avg_disc_cmd_valid             : in std_logic;
    l_avg_disc_cmd_ready             : out std_logic;
    l_avg_disc_cmd_firstIdx          : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    l_avg_disc_cmd_lastIdx           : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    l_avg_disc_cmd_ctrl              : in std_logic_vector(L_AVG_DISC_BUS_ADDR_WIDTH - 1 downto 0);
    l_avg_disc_cmd_tag               : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    l_avg_disc_unl_valid             : out std_logic;
    l_avg_disc_unl_ready             : in std_logic;
    l_avg_disc_unl_tag               : out std_logic_vector(TAG_WIDTH - 1 downto 0);
    l_count_order_valid              : in std_logic;
    l_count_order_ready              : out std_logic;
    l_count_order_dvalid             : in std_logic;
    l_count_order_last               : in std_logic;
    l_count_order                    : in std_logic_vector(63 downto 0);
    l_count_order_bus_wreq_valid     : out std_logic;
    l_count_order_bus_wreq_ready     : in std_logic;
    l_count_order_bus_wreq_addr      : out std_logic_vector(L_COUNT_ORDER_BUS_ADDR_WIDTH - 1 downto 0);
    l_count_order_bus_wreq_len       : out std_logic_vector(L_COUNT_ORDER_BUS_LEN_WIDTH - 1 downto 0);
    l_count_order_bus_wreq_last      : out std_logic;
    l_count_order_bus_wdat_valid     : out std_logic;
    l_count_order_bus_wdat_ready     : in std_logic;
    l_count_order_bus_wdat_data      : out std_logic_vector(L_COUNT_ORDER_BUS_DATA_WIDTH - 1 downto 0);
    l_count_order_bus_wdat_strobe    : out std_logic_vector(L_COUNT_ORDER_BUS_DATA_WIDTH/8 - 1 downto 0);
    l_count_order_bus_wdat_last      : out std_logic;
    l_count_order_bus_wrep_valid     : in std_logic;
    l_count_order_bus_wrep_ready     : out std_logic;
    l_count_order_bus_wrep_ok        : in std_logic;
    l_count_order_cmd_valid          : in std_logic;
    l_count_order_cmd_ready          : out std_logic;
    l_count_order_cmd_firstIdx       : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    l_count_order_cmd_lastIdx        : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
    l_count_order_cmd_ctrl           : in std_logic_vector(L_COUNT_ORDER_BUS_ADDR_WIDTH - 1 downto 0);
    l_count_order_cmd_tag            : in std_logic_vector(TAG_WIDTH - 1 downto 0);
    l_count_order_unl_valid          : out std_logic;
    l_count_order_unl_ready          : in std_logic;
    l_count_order_unl_tag            : out std_logic_vector(TAG_WIDTH - 1 downto 0)
  );
end entity;

architecture Implementation of PriceSummary_l is
  signal quantity_inst_cmd_valid             : std_logic;
  signal quantity_inst_cmd_ready             : std_logic;
  signal quantity_inst_cmd_firstIdx          : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal quantity_inst_cmd_lastIdx           : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal quantity_inst_cmd_ctrl              : std_logic_vector(L_QUANTITY_BUS_ADDR_WIDTH - 1 downto 0);
  signal quantity_inst_cmd_tag               : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal quantity_inst_unl_valid             : std_logic;
  signal quantity_inst_unl_ready             : std_logic;
  signal quantity_inst_unl_tag               : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal quantity_inst_bus_rreq_valid        : std_logic;
  signal quantity_inst_bus_rreq_ready        : std_logic;
  signal quantity_inst_bus_rreq_addr         : std_logic_vector(L_QUANTITY_BUS_ADDR_WIDTH - 1 downto 0);
  signal quantity_inst_bus_rreq_len          : std_logic_vector(L_QUANTITY_BUS_LEN_WIDTH - 1 downto 0);
  signal quantity_inst_bus_rdat_valid        : std_logic;
  signal quantity_inst_bus_rdat_ready        : std_logic;
  signal quantity_inst_bus_rdat_data         : std_logic_vector(L_QUANTITY_BUS_DATA_WIDTH - 1 downto 0);
  signal quantity_inst_bus_rdat_last         : std_logic;

  signal quantity_inst_out_valid             : std_logic_vector(0 downto 0);
  signal quantity_inst_out_ready             : std_logic_vector(0 downto 0);
  signal quantity_inst_out_data              : std_logic_vector(63 downto 0);
  signal quantity_inst_out_dvalid            : std_logic_vector(0 downto 0);
  signal quantity_inst_out_last              : std_logic_vector(0 downto 0);

  signal extendedprice_inst_cmd_valid        : std_logic;
  signal extendedprice_inst_cmd_ready        : std_logic;
  signal extendedprice_inst_cmd_firstIdx     : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal extendedprice_inst_cmd_lastIdx      : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal extendedprice_inst_cmd_ctrl         : std_logic_vector(L_EXTENDEDPRICE_BUS_ADDR_WIDTH - 1 downto 0);
  signal extendedprice_inst_cmd_tag          : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal extendedprice_inst_unl_valid        : std_logic;
  signal extendedprice_inst_unl_ready        : std_logic;
  signal extendedprice_inst_unl_tag          : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal extendedprice_inst_bus_rreq_valid   : std_logic;
  signal extendedprice_inst_bus_rreq_ready   : std_logic;
  signal extendedprice_inst_bus_rreq_addr    : std_logic_vector(L_EXTENDEDPRICE_BUS_ADDR_WIDTH - 1 downto 0);
  signal extendedprice_inst_bus_rreq_len     : std_logic_vector(L_EXTENDEDPRICE_BUS_LEN_WIDTH - 1 downto 0);
  signal extendedprice_inst_bus_rdat_valid   : std_logic;
  signal extendedprice_inst_bus_rdat_ready   : std_logic;
  signal extendedprice_inst_bus_rdat_data    : std_logic_vector(L_EXTENDEDPRICE_BUS_DATA_WIDTH - 1 downto 0);
  signal extendedprice_inst_bus_rdat_last    : std_logic;

  signal extendedprice_inst_out_valid        : std_logic_vector(0 downto 0);
  signal extendedprice_inst_out_ready        : std_logic_vector(0 downto 0);
  signal extendedprice_inst_out_data         : std_logic_vector(63 downto 0);
  signal extendedprice_inst_out_dvalid       : std_logic_vector(0 downto 0);
  signal extendedprice_inst_out_last         : std_logic_vector(0 downto 0);

  signal discount_inst_cmd_valid             : std_logic;
  signal discount_inst_cmd_ready             : std_logic;
  signal discount_inst_cmd_firstIdx          : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal discount_inst_cmd_lastIdx           : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal discount_inst_cmd_ctrl              : std_logic_vector(L_DISCOUNT_BUS_ADDR_WIDTH - 1 downto 0);
  signal discount_inst_cmd_tag               : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal discount_inst_unl_valid             : std_logic;
  signal discount_inst_unl_ready             : std_logic;
  signal discount_inst_unl_tag               : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal discount_inst_bus_rreq_valid        : std_logic;
  signal discount_inst_bus_rreq_ready        : std_logic;
  signal discount_inst_bus_rreq_addr         : std_logic_vector(L_DISCOUNT_BUS_ADDR_WIDTH - 1 downto 0);
  signal discount_inst_bus_rreq_len          : std_logic_vector(L_DISCOUNT_BUS_LEN_WIDTH - 1 downto 0);
  signal discount_inst_bus_rdat_valid        : std_logic;
  signal discount_inst_bus_rdat_ready        : std_logic;
  signal discount_inst_bus_rdat_data         : std_logic_vector(L_DISCOUNT_BUS_DATA_WIDTH - 1 downto 0);
  signal discount_inst_bus_rdat_last         : std_logic;

  signal discount_inst_out_valid             : std_logic_vector(0 downto 0);
  signal discount_inst_out_ready             : std_logic_vector(0 downto 0);
  signal discount_inst_out_data              : std_logic_vector(63 downto 0);
  signal discount_inst_out_dvalid            : std_logic_vector(0 downto 0);
  signal discount_inst_out_last              : std_logic_vector(0 downto 0);

  signal tax_inst_cmd_valid                  : std_logic;
  signal tax_inst_cmd_ready                  : std_logic;
  signal tax_inst_cmd_firstIdx               : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal tax_inst_cmd_lastIdx                : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal tax_inst_cmd_ctrl                   : std_logic_vector(L_TAX_BUS_ADDR_WIDTH - 1 downto 0);
  signal tax_inst_cmd_tag                    : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal tax_inst_unl_valid                  : std_logic;
  signal tax_inst_unl_ready                  : std_logic;
  signal tax_inst_unl_tag                    : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal tax_inst_bus_rreq_valid             : std_logic;
  signal tax_inst_bus_rreq_ready             : std_logic;
  signal tax_inst_bus_rreq_addr              : std_logic_vector(L_TAX_BUS_ADDR_WIDTH - 1 downto 0);
  signal tax_inst_bus_rreq_len               : std_logic_vector(L_TAX_BUS_LEN_WIDTH - 1 downto 0);
  signal tax_inst_bus_rdat_valid             : std_logic;
  signal tax_inst_bus_rdat_ready             : std_logic;
  signal tax_inst_bus_rdat_data              : std_logic_vector(L_TAX_BUS_DATA_WIDTH - 1 downto 0);
  signal tax_inst_bus_rdat_last              : std_logic;

  signal tax_inst_out_valid                  : std_logic_vector(0 downto 0);
  signal tax_inst_out_ready                  : std_logic_vector(0 downto 0);
  signal tax_inst_out_data                   : std_logic_vector(63 downto 0);
  signal tax_inst_out_dvalid                 : std_logic_vector(0 downto 0);
  signal tax_inst_out_last                   : std_logic_vector(0 downto 0);

  signal returnflag_inst_cmd_valid           : std_logic;
  signal returnflag_inst_cmd_ready           : std_logic;
  signal returnflag_inst_cmd_firstIdx        : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal returnflag_inst_cmd_lastIdx         : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal returnflag_inst_cmd_ctrl            : std_logic_vector(L_RETURNFLAG_BUS_ADDR_WIDTH * 2 - 1 downto 0);
  signal returnflag_inst_cmd_tag             : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal returnflag_inst_unl_valid           : std_logic;
  signal returnflag_inst_unl_ready           : std_logic;
  signal returnflag_inst_unl_tag             : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal returnflag_inst_bus_rreq_valid      : std_logic;
  signal returnflag_inst_bus_rreq_ready      : std_logic;
  signal returnflag_inst_bus_rreq_addr       : std_logic_vector(L_RETURNFLAG_BUS_ADDR_WIDTH - 1 downto 0);
  signal returnflag_inst_bus_rreq_len        : std_logic_vector(L_RETURNFLAG_BUS_LEN_WIDTH - 1 downto 0);
  signal returnflag_inst_bus_rdat_valid      : std_logic;
  signal returnflag_inst_bus_rdat_ready      : std_logic;
  signal returnflag_inst_bus_rdat_data       : std_logic_vector(L_RETURNFLAG_BUS_DATA_WIDTH - 1 downto 0);
  signal returnflag_inst_bus_rdat_last       : std_logic;

  signal returnflag_inst_out_valid           : std_logic_vector(1 downto 0);
  signal returnflag_inst_out_ready           : std_logic_vector(1 downto 0);
  signal returnflag_inst_out_data            : std_logic_vector(41 downto 0);
  signal returnflag_inst_out_dvalid          : std_logic_vector(1 downto 0);
  signal returnflag_inst_out_last            : std_logic_vector(1 downto 0);

  signal linestatus_inst_cmd_valid           : std_logic;
  signal linestatus_inst_cmd_ready           : std_logic;
  signal linestatus_inst_cmd_firstIdx        : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal linestatus_inst_cmd_lastIdx         : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal linestatus_inst_cmd_ctrl            : std_logic_vector(L_LINESTATUS_BUS_ADDR_WIDTH * 2 - 1 downto 0);
  signal linestatus_inst_cmd_tag             : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal linestatus_inst_unl_valid           : std_logic;
  signal linestatus_inst_unl_ready           : std_logic;
  signal linestatus_inst_unl_tag             : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal linestatus_inst_bus_rreq_valid      : std_logic;
  signal linestatus_inst_bus_rreq_ready      : std_logic;
  signal linestatus_inst_bus_rreq_addr       : std_logic_vector(L_LINESTATUS_BUS_ADDR_WIDTH - 1 downto 0);
  signal linestatus_inst_bus_rreq_len        : std_logic_vector(L_LINESTATUS_BUS_LEN_WIDTH - 1 downto 0);
  signal linestatus_inst_bus_rdat_valid      : std_logic;
  signal linestatus_inst_bus_rdat_ready      : std_logic;
  signal linestatus_inst_bus_rdat_data       : std_logic_vector(L_LINESTATUS_BUS_DATA_WIDTH - 1 downto 0);
  signal linestatus_inst_bus_rdat_last       : std_logic;

  signal linestatus_inst_out_valid           : std_logic_vector(1 downto 0);
  signal linestatus_inst_out_ready           : std_logic_vector(1 downto 0);
  signal linestatus_inst_out_data            : std_logic_vector(41 downto 0);
  signal linestatus_inst_out_dvalid          : std_logic_vector(1 downto 0);
  signal linestatus_inst_out_last            : std_logic_vector(1 downto 0);

  signal shipdate_inst_cmd_valid             : std_logic;
  signal shipdate_inst_cmd_ready             : std_logic;
  signal shipdate_inst_cmd_firstIdx          : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal shipdate_inst_cmd_lastIdx           : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal shipdate_inst_cmd_ctrl              : std_logic_vector(L_SHIPDATE_BUS_ADDR_WIDTH - 1 downto 0);
  signal shipdate_inst_cmd_tag               : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal shipdate_inst_unl_valid             : std_logic;
  signal shipdate_inst_unl_ready             : std_logic;
  signal shipdate_inst_unl_tag               : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal shipdate_inst_bus_rreq_valid        : std_logic;
  signal shipdate_inst_bus_rreq_ready        : std_logic;
  signal shipdate_inst_bus_rreq_addr         : std_logic_vector(L_SHIPDATE_BUS_ADDR_WIDTH - 1 downto 0);
  signal shipdate_inst_bus_rreq_len          : std_logic_vector(L_SHIPDATE_BUS_LEN_WIDTH - 1 downto 0);
  signal shipdate_inst_bus_rdat_valid        : std_logic;
  signal shipdate_inst_bus_rdat_ready        : std_logic;
  signal shipdate_inst_bus_rdat_data         : std_logic_vector(L_SHIPDATE_BUS_DATA_WIDTH - 1 downto 0);
  signal shipdate_inst_bus_rdat_last         : std_logic;

  signal shipdate_inst_out_valid             : std_logic_vector(0 downto 0);
  signal shipdate_inst_out_ready             : std_logic_vector(0 downto 0);
  signal shipdate_inst_out_data              : std_logic_vector(31 downto 0);
  signal shipdate_inst_out_dvalid            : std_logic_vector(0 downto 0);
  signal shipdate_inst_out_last              : std_logic_vector(0 downto 0);

  signal returnflag_o_inst_cmd_valid         : std_logic;
  signal returnflag_o_inst_cmd_ready         : std_logic;
  signal returnflag_o_inst_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal returnflag_o_inst_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal returnflag_o_inst_cmd_ctrl          : std_logic_vector(L_RETURNFLAG_O_BUS_ADDR_WIDTH * 2 - 1 downto 0);
  signal returnflag_o_inst_cmd_tag           : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal returnflag_o_inst_unl_valid         : std_logic;
  signal returnflag_o_inst_unl_ready         : std_logic;
  signal returnflag_o_inst_unl_tag           : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal returnflag_o_inst_bus_wreq_valid    : std_logic;
  signal returnflag_o_inst_bus_wreq_ready    : std_logic;
  signal returnflag_o_inst_bus_wreq_addr     : std_logic_vector(L_RETURNFLAG_O_BUS_ADDR_WIDTH - 1 downto 0);
  signal returnflag_o_inst_bus_wreq_len      : std_logic_vector(L_RETURNFLAG_O_BUS_LEN_WIDTH - 1 downto 0);
  signal returnflag_o_inst_bus_wreq_last     : std_logic;
  signal returnflag_o_inst_bus_wdat_valid    : std_logic;
  signal returnflag_o_inst_bus_wdat_ready    : std_logic;
  signal returnflag_o_inst_bus_wdat_data     : std_logic_vector(L_RETURNFLAG_O_BUS_DATA_WIDTH - 1 downto 0);
  signal returnflag_o_inst_bus_wdat_strobe   : std_logic_vector(L_RETURNFLAG_O_BUS_DATA_WIDTH/8 - 1 downto 0);
  signal returnflag_o_inst_bus_wdat_last     : std_logic;
  signal returnflag_o_inst_bus_wrep_valid    : std_logic;
  signal returnflag_o_inst_bus_wrep_ready    : std_logic;
  signal returnflag_o_inst_bus_wrep_ok       : std_logic;

  signal returnflag_o_inst_in_valid          : std_logic_vector(1 downto 0);
  signal returnflag_o_inst_in_ready          : std_logic_vector(1 downto 0);
  signal returnflag_o_inst_in_data           : std_logic_vector(41 downto 0);
  signal returnflag_o_inst_in_dvalid         : std_logic_vector(1 downto 0);
  signal returnflag_o_inst_in_last           : std_logic_vector(1 downto 0);

  signal linestatus_o_inst_cmd_valid         : std_logic;
  signal linestatus_o_inst_cmd_ready         : std_logic;
  signal linestatus_o_inst_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal linestatus_o_inst_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal linestatus_o_inst_cmd_ctrl          : std_logic_vector(L_LINESTATUS_O_BUS_ADDR_WIDTH * 2 - 1 downto 0);
  signal linestatus_o_inst_cmd_tag           : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal linestatus_o_inst_unl_valid         : std_logic;
  signal linestatus_o_inst_unl_ready         : std_logic;
  signal linestatus_o_inst_unl_tag           : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal linestatus_o_inst_bus_wreq_valid    : std_logic;
  signal linestatus_o_inst_bus_wreq_ready    : std_logic;
  signal linestatus_o_inst_bus_wreq_addr     : std_logic_vector(L_LINESTATUS_O_BUS_ADDR_WIDTH - 1 downto 0);
  signal linestatus_o_inst_bus_wreq_len      : std_logic_vector(L_LINESTATUS_O_BUS_LEN_WIDTH - 1 downto 0);
  signal linestatus_o_inst_bus_wreq_last     : std_logic;
  signal linestatus_o_inst_bus_wdat_valid    : std_logic;
  signal linestatus_o_inst_bus_wdat_ready    : std_logic;
  signal linestatus_o_inst_bus_wdat_data     : std_logic_vector(L_LINESTATUS_O_BUS_DATA_WIDTH - 1 downto 0);
  signal linestatus_o_inst_bus_wdat_strobe   : std_logic_vector(L_LINESTATUS_O_BUS_DATA_WIDTH/8 - 1 downto 0);
  signal linestatus_o_inst_bus_wdat_last     : std_logic;
  signal linestatus_o_inst_bus_wrep_valid    : std_logic;
  signal linestatus_o_inst_bus_wrep_ready    : std_logic;
  signal linestatus_o_inst_bus_wrep_ok       : std_logic;

  signal linestatus_o_inst_in_valid          : std_logic_vector(1 downto 0);
  signal linestatus_o_inst_in_ready          : std_logic_vector(1 downto 0);
  signal linestatus_o_inst_in_data           : std_logic_vector(41 downto 0);
  signal linestatus_o_inst_in_dvalid         : std_logic_vector(1 downto 0);
  signal linestatus_o_inst_in_last           : std_logic_vector(1 downto 0);

  signal sum_qty_inst_cmd_valid              : std_logic;
  signal sum_qty_inst_cmd_ready              : std_logic;
  signal sum_qty_inst_cmd_firstIdx           : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal sum_qty_inst_cmd_lastIdx            : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal sum_qty_inst_cmd_ctrl               : std_logic_vector(L_SUM_QTY_BUS_ADDR_WIDTH - 1 downto 0);
  signal sum_qty_inst_cmd_tag                : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal sum_qty_inst_unl_valid              : std_logic;
  signal sum_qty_inst_unl_ready              : std_logic;
  signal sum_qty_inst_unl_tag                : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal sum_qty_inst_bus_wreq_valid         : std_logic;
  signal sum_qty_inst_bus_wreq_ready         : std_logic;
  signal sum_qty_inst_bus_wreq_addr          : std_logic_vector(L_SUM_QTY_BUS_ADDR_WIDTH - 1 downto 0);
  signal sum_qty_inst_bus_wreq_len           : std_logic_vector(L_SUM_QTY_BUS_LEN_WIDTH - 1 downto 0);
  signal sum_qty_inst_bus_wreq_last          : std_logic;
  signal sum_qty_inst_bus_wdat_valid         : std_logic;
  signal sum_qty_inst_bus_wdat_ready         : std_logic;
  signal sum_qty_inst_bus_wdat_data          : std_logic_vector(L_SUM_QTY_BUS_DATA_WIDTH - 1 downto 0);
  signal sum_qty_inst_bus_wdat_strobe        : std_logic_vector(L_SUM_QTY_BUS_DATA_WIDTH/8 - 1 downto 0);
  signal sum_qty_inst_bus_wdat_last          : std_logic;
  signal sum_qty_inst_bus_wrep_valid         : std_logic;
  signal sum_qty_inst_bus_wrep_ready         : std_logic;
  signal sum_qty_inst_bus_wrep_ok            : std_logic;

  signal sum_qty_inst_in_valid               : std_logic_vector(0 downto 0);
  signal sum_qty_inst_in_ready               : std_logic_vector(0 downto 0);
  signal sum_qty_inst_in_data                : std_logic_vector(63 downto 0);
  signal sum_qty_inst_in_dvalid              : std_logic_vector(0 downto 0);
  signal sum_qty_inst_in_last                : std_logic_vector(0 downto 0);

  signal sum_base_price_inst_cmd_valid       : std_logic;
  signal sum_base_price_inst_cmd_ready       : std_logic;
  signal sum_base_price_inst_cmd_firstIdx    : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal sum_base_price_inst_cmd_lastIdx     : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal sum_base_price_inst_cmd_ctrl        : std_logic_vector(L_SUM_BASE_PRICE_BUS_ADDR_WIDTH - 1 downto 0);
  signal sum_base_price_inst_cmd_tag         : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal sum_base_price_inst_unl_valid       : std_logic;
  signal sum_base_price_inst_unl_ready       : std_logic;
  signal sum_base_price_inst_unl_tag         : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal sum_base_price_inst_bus_wreq_valid  : std_logic;
  signal sum_base_price_inst_bus_wreq_ready  : std_logic;
  signal sum_base_price_inst_bus_wreq_addr   : std_logic_vector(L_SUM_BASE_PRICE_BUS_ADDR_WIDTH - 1 downto 0);
  signal sum_base_price_inst_bus_wreq_len    : std_logic_vector(L_SUM_BASE_PRICE_BUS_LEN_WIDTH - 1 downto 0);
  signal sum_base_price_inst_bus_wreq_last   : std_logic;
  signal sum_base_price_inst_bus_wdat_valid  : std_logic;
  signal sum_base_price_inst_bus_wdat_ready  : std_logic;
  signal sum_base_price_inst_bus_wdat_data   : std_logic_vector(L_SUM_BASE_PRICE_BUS_DATA_WIDTH - 1 downto 0);
  signal sum_base_price_inst_bus_wdat_strobe : std_logic_vector(L_SUM_BASE_PRICE_BUS_DATA_WIDTH/8 - 1 downto 0);
  signal sum_base_price_inst_bus_wdat_last   : std_logic;
  signal sum_base_price_inst_bus_wrep_valid  : std_logic;
  signal sum_base_price_inst_bus_wrep_ready  : std_logic;
  signal sum_base_price_inst_bus_wrep_ok     : std_logic;

  signal sum_base_price_inst_in_valid        : std_logic_vector(0 downto 0);
  signal sum_base_price_inst_in_ready        : std_logic_vector(0 downto 0);
  signal sum_base_price_inst_in_data         : std_logic_vector(63 downto 0);
  signal sum_base_price_inst_in_dvalid       : std_logic_vector(0 downto 0);
  signal sum_base_price_inst_in_last         : std_logic_vector(0 downto 0);

  signal sum_disc_price_inst_cmd_valid       : std_logic;
  signal sum_disc_price_inst_cmd_ready       : std_logic;
  signal sum_disc_price_inst_cmd_firstIdx    : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal sum_disc_price_inst_cmd_lastIdx     : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal sum_disc_price_inst_cmd_ctrl        : std_logic_vector(L_SUM_DISC_PRICE_BUS_ADDR_WIDTH - 1 downto 0);
  signal sum_disc_price_inst_cmd_tag         : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal sum_disc_price_inst_unl_valid       : std_logic;
  signal sum_disc_price_inst_unl_ready       : std_logic;
  signal sum_disc_price_inst_unl_tag         : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal sum_disc_price_inst_bus_wreq_valid  : std_logic;
  signal sum_disc_price_inst_bus_wreq_ready  : std_logic;
  signal sum_disc_price_inst_bus_wreq_addr   : std_logic_vector(L_SUM_DISC_PRICE_BUS_ADDR_WIDTH - 1 downto 0);
  signal sum_disc_price_inst_bus_wreq_len    : std_logic_vector(L_SUM_DISC_PRICE_BUS_LEN_WIDTH - 1 downto 0);
  signal sum_disc_price_inst_bus_wreq_last   : std_logic;
  signal sum_disc_price_inst_bus_wdat_valid  : std_logic;
  signal sum_disc_price_inst_bus_wdat_ready  : std_logic;
  signal sum_disc_price_inst_bus_wdat_data   : std_logic_vector(L_SUM_DISC_PRICE_BUS_DATA_WIDTH - 1 downto 0);
  signal sum_disc_price_inst_bus_wdat_strobe : std_logic_vector(L_SUM_DISC_PRICE_BUS_DATA_WIDTH/8 - 1 downto 0);
  signal sum_disc_price_inst_bus_wdat_last   : std_logic;
  signal sum_disc_price_inst_bus_wrep_valid  : std_logic;
  signal sum_disc_price_inst_bus_wrep_ready  : std_logic;
  signal sum_disc_price_inst_bus_wrep_ok     : std_logic;

  signal sum_disc_price_inst_in_valid        : std_logic_vector(0 downto 0);
  signal sum_disc_price_inst_in_ready        : std_logic_vector(0 downto 0);
  signal sum_disc_price_inst_in_data         : std_logic_vector(63 downto 0);
  signal sum_disc_price_inst_in_dvalid       : std_logic_vector(0 downto 0);
  signal sum_disc_price_inst_in_last         : std_logic_vector(0 downto 0);

  signal sum_charge_inst_cmd_valid           : std_logic;
  signal sum_charge_inst_cmd_ready           : std_logic;
  signal sum_charge_inst_cmd_firstIdx        : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal sum_charge_inst_cmd_lastIdx         : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal sum_charge_inst_cmd_ctrl            : std_logic_vector(L_SUM_CHARGE_BUS_ADDR_WIDTH - 1 downto 0);
  signal sum_charge_inst_cmd_tag             : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal sum_charge_inst_unl_valid           : std_logic;
  signal sum_charge_inst_unl_ready           : std_logic;
  signal sum_charge_inst_unl_tag             : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal sum_charge_inst_bus_wreq_valid      : std_logic;
  signal sum_charge_inst_bus_wreq_ready      : std_logic;
  signal sum_charge_inst_bus_wreq_addr       : std_logic_vector(L_SUM_CHARGE_BUS_ADDR_WIDTH - 1 downto 0);
  signal sum_charge_inst_bus_wreq_len        : std_logic_vector(L_SUM_CHARGE_BUS_LEN_WIDTH - 1 downto 0);
  signal sum_charge_inst_bus_wreq_last       : std_logic;
  signal sum_charge_inst_bus_wdat_valid      : std_logic;
  signal sum_charge_inst_bus_wdat_ready      : std_logic;
  signal sum_charge_inst_bus_wdat_data       : std_logic_vector(L_SUM_CHARGE_BUS_DATA_WIDTH - 1 downto 0);
  signal sum_charge_inst_bus_wdat_strobe     : std_logic_vector(L_SUM_CHARGE_BUS_DATA_WIDTH/8 - 1 downto 0);
  signal sum_charge_inst_bus_wdat_last       : std_logic;
  signal sum_charge_inst_bus_wrep_valid      : std_logic;
  signal sum_charge_inst_bus_wrep_ready      : std_logic;
  signal sum_charge_inst_bus_wrep_ok         : std_logic;

  signal sum_charge_inst_in_valid            : std_logic_vector(0 downto 0);
  signal sum_charge_inst_in_ready            : std_logic_vector(0 downto 0);
  signal sum_charge_inst_in_data             : std_logic_vector(63 downto 0);
  signal sum_charge_inst_in_dvalid           : std_logic_vector(0 downto 0);
  signal sum_charge_inst_in_last             : std_logic_vector(0 downto 0);

  signal avg_qty_inst_cmd_valid              : std_logic;
  signal avg_qty_inst_cmd_ready              : std_logic;
  signal avg_qty_inst_cmd_firstIdx           : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal avg_qty_inst_cmd_lastIdx            : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal avg_qty_inst_cmd_ctrl               : std_logic_vector(L_AVG_QTY_BUS_ADDR_WIDTH - 1 downto 0);
  signal avg_qty_inst_cmd_tag                : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal avg_qty_inst_unl_valid              : std_logic;
  signal avg_qty_inst_unl_ready              : std_logic;
  signal avg_qty_inst_unl_tag                : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal avg_qty_inst_bus_wreq_valid         : std_logic;
  signal avg_qty_inst_bus_wreq_ready         : std_logic;
  signal avg_qty_inst_bus_wreq_addr          : std_logic_vector(L_AVG_QTY_BUS_ADDR_WIDTH - 1 downto 0);
  signal avg_qty_inst_bus_wreq_len           : std_logic_vector(L_AVG_QTY_BUS_LEN_WIDTH - 1 downto 0);
  signal avg_qty_inst_bus_wreq_last          : std_logic;
  signal avg_qty_inst_bus_wdat_valid         : std_logic;
  signal avg_qty_inst_bus_wdat_ready         : std_logic;
  signal avg_qty_inst_bus_wdat_data          : std_logic_vector(L_AVG_QTY_BUS_DATA_WIDTH - 1 downto 0);
  signal avg_qty_inst_bus_wdat_strobe        : std_logic_vector(L_AVG_QTY_BUS_DATA_WIDTH/8 - 1 downto 0);
  signal avg_qty_inst_bus_wdat_last          : std_logic;
  signal avg_qty_inst_bus_wrep_valid         : std_logic;
  signal avg_qty_inst_bus_wrep_ready         : std_logic;
  signal avg_qty_inst_bus_wrep_ok            : std_logic;

  signal avg_qty_inst_in_valid               : std_logic_vector(0 downto 0);
  signal avg_qty_inst_in_ready               : std_logic_vector(0 downto 0);
  signal avg_qty_inst_in_data                : std_logic_vector(63 downto 0);
  signal avg_qty_inst_in_dvalid              : std_logic_vector(0 downto 0);
  signal avg_qty_inst_in_last                : std_logic_vector(0 downto 0);

  signal avg_price_inst_cmd_valid            : std_logic;
  signal avg_price_inst_cmd_ready            : std_logic;
  signal avg_price_inst_cmd_firstIdx         : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal avg_price_inst_cmd_lastIdx          : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal avg_price_inst_cmd_ctrl             : std_logic_vector(L_AVG_PRICE_BUS_ADDR_WIDTH - 1 downto 0);
  signal avg_price_inst_cmd_tag              : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal avg_price_inst_unl_valid            : std_logic;
  signal avg_price_inst_unl_ready            : std_logic;
  signal avg_price_inst_unl_tag              : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal avg_price_inst_bus_wreq_valid       : std_logic;
  signal avg_price_inst_bus_wreq_ready       : std_logic;
  signal avg_price_inst_bus_wreq_addr        : std_logic_vector(L_AVG_PRICE_BUS_ADDR_WIDTH - 1 downto 0);
  signal avg_price_inst_bus_wreq_len         : std_logic_vector(L_AVG_PRICE_BUS_LEN_WIDTH - 1 downto 0);
  signal avg_price_inst_bus_wreq_last        : std_logic;
  signal avg_price_inst_bus_wdat_valid       : std_logic;
  signal avg_price_inst_bus_wdat_ready       : std_logic;
  signal avg_price_inst_bus_wdat_data        : std_logic_vector(L_AVG_PRICE_BUS_DATA_WIDTH - 1 downto 0);
  signal avg_price_inst_bus_wdat_strobe      : std_logic_vector(L_AVG_PRICE_BUS_DATA_WIDTH/8 - 1 downto 0);
  signal avg_price_inst_bus_wdat_last        : std_logic;
  signal avg_price_inst_bus_wrep_valid       : std_logic;
  signal avg_price_inst_bus_wrep_ready       : std_logic;
  signal avg_price_inst_bus_wrep_ok          : std_logic;

  signal avg_price_inst_in_valid             : std_logic_vector(0 downto 0);
  signal avg_price_inst_in_ready             : std_logic_vector(0 downto 0);
  signal avg_price_inst_in_data              : std_logic_vector(63 downto 0);
  signal avg_price_inst_in_dvalid            : std_logic_vector(0 downto 0);
  signal avg_price_inst_in_last              : std_logic_vector(0 downto 0);

  signal avg_disc_inst_cmd_valid             : std_logic;
  signal avg_disc_inst_cmd_ready             : std_logic;
  signal avg_disc_inst_cmd_firstIdx          : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal avg_disc_inst_cmd_lastIdx           : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal avg_disc_inst_cmd_ctrl              : std_logic_vector(L_AVG_DISC_BUS_ADDR_WIDTH - 1 downto 0);
  signal avg_disc_inst_cmd_tag               : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal avg_disc_inst_unl_valid             : std_logic;
  signal avg_disc_inst_unl_ready             : std_logic;
  signal avg_disc_inst_unl_tag               : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal avg_disc_inst_bus_wreq_valid        : std_logic;
  signal avg_disc_inst_bus_wreq_ready        : std_logic;
  signal avg_disc_inst_bus_wreq_addr         : std_logic_vector(L_AVG_DISC_BUS_ADDR_WIDTH - 1 downto 0);
  signal avg_disc_inst_bus_wreq_len          : std_logic_vector(L_AVG_DISC_BUS_LEN_WIDTH - 1 downto 0);
  signal avg_disc_inst_bus_wreq_last         : std_logic;
  signal avg_disc_inst_bus_wdat_valid        : std_logic;
  signal avg_disc_inst_bus_wdat_ready        : std_logic;
  signal avg_disc_inst_bus_wdat_data         : std_logic_vector(L_AVG_DISC_BUS_DATA_WIDTH - 1 downto 0);
  signal avg_disc_inst_bus_wdat_strobe       : std_logic_vector(L_AVG_DISC_BUS_DATA_WIDTH/8 - 1 downto 0);
  signal avg_disc_inst_bus_wdat_last         : std_logic;
  signal avg_disc_inst_bus_wrep_valid        : std_logic;
  signal avg_disc_inst_bus_wrep_ready        : std_logic;
  signal avg_disc_inst_bus_wrep_ok           : std_logic;

  signal avg_disc_inst_in_valid              : std_logic_vector(0 downto 0);
  signal avg_disc_inst_in_ready              : std_logic_vector(0 downto 0);
  signal avg_disc_inst_in_data               : std_logic_vector(63 downto 0);
  signal avg_disc_inst_in_dvalid             : std_logic_vector(0 downto 0);
  signal avg_disc_inst_in_last               : std_logic_vector(0 downto 0);

  signal count_order_inst_cmd_valid          : std_logic;
  signal count_order_inst_cmd_ready          : std_logic;
  signal count_order_inst_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal count_order_inst_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal count_order_inst_cmd_ctrl           : std_logic_vector(L_COUNT_ORDER_BUS_ADDR_WIDTH - 1 downto 0);
  signal count_order_inst_cmd_tag            : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal count_order_inst_unl_valid          : std_logic;
  signal count_order_inst_unl_ready          : std_logic;
  signal count_order_inst_unl_tag            : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal count_order_inst_bus_wreq_valid     : std_logic;
  signal count_order_inst_bus_wreq_ready     : std_logic;
  signal count_order_inst_bus_wreq_addr      : std_logic_vector(L_COUNT_ORDER_BUS_ADDR_WIDTH - 1 downto 0);
  signal count_order_inst_bus_wreq_len       : std_logic_vector(L_COUNT_ORDER_BUS_LEN_WIDTH - 1 downto 0);
  signal count_order_inst_bus_wreq_last      : std_logic;
  signal count_order_inst_bus_wdat_valid     : std_logic;
  signal count_order_inst_bus_wdat_ready     : std_logic;
  signal count_order_inst_bus_wdat_data      : std_logic_vector(L_COUNT_ORDER_BUS_DATA_WIDTH - 1 downto 0);
  signal count_order_inst_bus_wdat_strobe    : std_logic_vector(L_COUNT_ORDER_BUS_DATA_WIDTH/8 - 1 downto 0);
  signal count_order_inst_bus_wdat_last      : std_logic;
  signal count_order_inst_bus_wrep_valid     : std_logic;
  signal count_order_inst_bus_wrep_ready     : std_logic;
  signal count_order_inst_bus_wrep_ok        : std_logic;

  signal count_order_inst_in_valid           : std_logic_vector(0 downto 0);
  signal count_order_inst_in_ready           : std_logic_vector(0 downto 0);
  signal count_order_inst_in_data            : std_logic_vector(63 downto 0);
  signal count_order_inst_in_dvalid          : std_logic_vector(0 downto 0);
  signal count_order_inst_in_last            : std_logic_vector(0 downto 0);

begin
  returnflag_o_inst : ArrayWriter
  generic map(
    BUS_ADDR_WIDTH     => L_RETURNFLAG_O_BUS_ADDR_WIDTH,
    BUS_DATA_WIDTH     => L_RETURNFLAG_O_BUS_DATA_WIDTH,
    BUS_LEN_WIDTH      => L_RETURNFLAG_O_BUS_LEN_WIDTH,
    BUS_BURST_STEP_LEN => L_RETURNFLAG_O_BUS_BURST_STEP_LEN,
    BUS_BURST_MAX_LEN  => L_RETURNFLAG_O_BUS_BURST_MAX_LEN,
    INDEX_WIDTH        => INDEX_WIDTH,
    CFG                => "listprim(8)",
    CMD_TAG_ENABLE     => true,
    CMD_TAG_WIDTH      => TAG_WIDTH
  )
  port map(
    bcd_clk         => bcd_clk,
    bcd_reset       => bcd_reset,
    kcd_clk         => kcd_clk,
    kcd_reset       => kcd_reset,
    cmd_valid       => returnflag_o_inst_cmd_valid,
    cmd_ready       => returnflag_o_inst_cmd_ready,
    cmd_firstIdx    => returnflag_o_inst_cmd_firstIdx,
    cmd_lastIdx     => returnflag_o_inst_cmd_lastIdx,
    cmd_ctrl        => returnflag_o_inst_cmd_ctrl,
    cmd_tag         => returnflag_o_inst_cmd_tag,
    unl_valid       => returnflag_o_inst_unl_valid,
    unl_ready       => returnflag_o_inst_unl_ready,
    unl_tag         => returnflag_o_inst_unl_tag,
    bus_wreq_valid  => returnflag_o_inst_bus_wreq_valid,
    bus_wreq_ready  => returnflag_o_inst_bus_wreq_ready,
    bus_wreq_addr   => returnflag_o_inst_bus_wreq_addr,
    bus_wreq_len    => returnflag_o_inst_bus_wreq_len,
    bus_wreq_last   => returnflag_o_inst_bus_wreq_last,
    bus_wdat_valid  => returnflag_o_inst_bus_wdat_valid,
    bus_wdat_ready  => returnflag_o_inst_bus_wdat_ready,
    bus_wdat_data   => returnflag_o_inst_bus_wdat_data,
    bus_wdat_strobe => returnflag_o_inst_bus_wdat_strobe,
    bus_wdat_last   => returnflag_o_inst_bus_wdat_last,
    bus_wrep_valid  => returnflag_o_inst_bus_wrep_valid,
    bus_wrep_ready  => returnflag_o_inst_bus_wrep_ready,
    bus_wrep_ok     => returnflag_o_inst_bus_wrep_ok,
    in_valid        => returnflag_o_inst_in_valid,
    in_ready        => returnflag_o_inst_in_ready,
    in_data         => returnflag_o_inst_in_data,
    in_dvalid       => returnflag_o_inst_in_dvalid,
    in_last         => returnflag_o_inst_in_last
  );

  linestatus_o_inst : ArrayWriter
  generic map(
    BUS_ADDR_WIDTH     => L_LINESTATUS_O_BUS_ADDR_WIDTH,
    BUS_DATA_WIDTH     => L_LINESTATUS_O_BUS_DATA_WIDTH,
    BUS_LEN_WIDTH      => L_LINESTATUS_O_BUS_LEN_WIDTH,
    BUS_BURST_STEP_LEN => L_LINESTATUS_O_BUS_BURST_STEP_LEN,
    BUS_BURST_MAX_LEN  => L_LINESTATUS_O_BUS_BURST_MAX_LEN,
    INDEX_WIDTH        => INDEX_WIDTH,
    CFG                => "listprim(8)",
    CMD_TAG_ENABLE     => true,
    CMD_TAG_WIDTH      => TAG_WIDTH
  )
  port map(
    bcd_clk         => bcd_clk,
    bcd_reset       => bcd_reset,
    kcd_clk         => kcd_clk,
    kcd_reset       => kcd_reset,
    cmd_valid       => linestatus_o_inst_cmd_valid,
    cmd_ready       => linestatus_o_inst_cmd_ready,
    cmd_firstIdx    => linestatus_o_inst_cmd_firstIdx,
    cmd_lastIdx     => linestatus_o_inst_cmd_lastIdx,
    cmd_ctrl        => linestatus_o_inst_cmd_ctrl,
    cmd_tag         => linestatus_o_inst_cmd_tag,
    unl_valid       => linestatus_o_inst_unl_valid,
    unl_ready       => linestatus_o_inst_unl_ready,
    unl_tag         => linestatus_o_inst_unl_tag,
    bus_wreq_valid  => linestatus_o_inst_bus_wreq_valid,
    bus_wreq_ready  => linestatus_o_inst_bus_wreq_ready,
    bus_wreq_addr   => linestatus_o_inst_bus_wreq_addr,
    bus_wreq_len    => linestatus_o_inst_bus_wreq_len,
    bus_wreq_last   => linestatus_o_inst_bus_wreq_last,
    bus_wdat_valid  => linestatus_o_inst_bus_wdat_valid,
    bus_wdat_ready  => linestatus_o_inst_bus_wdat_ready,
    bus_wdat_data   => linestatus_o_inst_bus_wdat_data,
    bus_wdat_strobe => linestatus_o_inst_bus_wdat_strobe,
    bus_wdat_last   => linestatus_o_inst_bus_wdat_last,
    bus_wrep_valid  => linestatus_o_inst_bus_wrep_valid,
    bus_wrep_ready  => linestatus_o_inst_bus_wrep_ready,
    bus_wrep_ok     => linestatus_o_inst_bus_wrep_ok,
    in_valid        => linestatus_o_inst_in_valid,
    in_ready        => linestatus_o_inst_in_ready,
    in_data         => linestatus_o_inst_in_data,
    in_dvalid       => linestatus_o_inst_in_dvalid,
    in_last         => linestatus_o_inst_in_last
  );

  sum_qty_inst : ArrayWriter
  generic map(
    BUS_ADDR_WIDTH     => L_SUM_QTY_BUS_ADDR_WIDTH,
    BUS_DATA_WIDTH     => L_SUM_QTY_BUS_DATA_WIDTH,
    BUS_LEN_WIDTH      => L_SUM_QTY_BUS_LEN_WIDTH,
    BUS_BURST_STEP_LEN => L_SUM_QTY_BUS_BURST_STEP_LEN,
    BUS_BURST_MAX_LEN  => L_SUM_QTY_BUS_BURST_MAX_LEN,
    INDEX_WIDTH        => INDEX_WIDTH,
    CFG                => "prim(64)",
    CMD_TAG_ENABLE     => true,
    CMD_TAG_WIDTH      => TAG_WIDTH
  )
  port map(
    bcd_clk         => bcd_clk,
    bcd_reset       => bcd_reset,
    kcd_clk         => kcd_clk,
    kcd_reset       => kcd_reset,
    cmd_valid       => sum_qty_inst_cmd_valid,
    cmd_ready       => sum_qty_inst_cmd_ready,
    cmd_firstIdx    => sum_qty_inst_cmd_firstIdx,
    cmd_lastIdx     => sum_qty_inst_cmd_lastIdx,
    cmd_ctrl        => sum_qty_inst_cmd_ctrl,
    cmd_tag         => sum_qty_inst_cmd_tag,
    unl_valid       => sum_qty_inst_unl_valid,
    unl_ready       => sum_qty_inst_unl_ready,
    unl_tag         => sum_qty_inst_unl_tag,
    bus_wreq_valid  => sum_qty_inst_bus_wreq_valid,
    bus_wreq_ready  => sum_qty_inst_bus_wreq_ready,
    bus_wreq_addr   => sum_qty_inst_bus_wreq_addr,
    bus_wreq_len    => sum_qty_inst_bus_wreq_len,
    bus_wreq_last   => sum_qty_inst_bus_wreq_last,
    bus_wdat_valid  => sum_qty_inst_bus_wdat_valid,
    bus_wdat_ready  => sum_qty_inst_bus_wdat_ready,
    bus_wdat_data   => sum_qty_inst_bus_wdat_data,
    bus_wdat_strobe => sum_qty_inst_bus_wdat_strobe,
    bus_wdat_last   => sum_qty_inst_bus_wdat_last,
    bus_wrep_valid  => sum_qty_inst_bus_wrep_valid,
    bus_wrep_ready  => sum_qty_inst_bus_wrep_ready,
    bus_wrep_ok     => sum_qty_inst_bus_wrep_ok,
    in_valid        => sum_qty_inst_in_valid,
    in_ready        => sum_qty_inst_in_ready,
    in_data         => sum_qty_inst_in_data,
    in_dvalid       => sum_qty_inst_in_dvalid,
    in_last         => sum_qty_inst_in_last
  );

  sum_base_price_inst : ArrayWriter
  generic map(
    BUS_ADDR_WIDTH     => L_SUM_BASE_PRICE_BUS_ADDR_WIDTH,
    BUS_DATA_WIDTH     => L_SUM_BASE_PRICE_BUS_DATA_WIDTH,
    BUS_LEN_WIDTH      => L_SUM_BASE_PRICE_BUS_LEN_WIDTH,
    BUS_BURST_STEP_LEN => L_SUM_BASE_PRICE_BUS_BURST_STEP_LEN,
    BUS_BURST_MAX_LEN  => L_SUM_BASE_PRICE_BUS_BURST_MAX_LEN,
    INDEX_WIDTH        => INDEX_WIDTH,
    CFG                => "prim(64)",
    CMD_TAG_ENABLE     => true,
    CMD_TAG_WIDTH      => TAG_WIDTH
  )
  port map(
    bcd_clk         => bcd_clk,
    bcd_reset       => bcd_reset,
    kcd_clk         => kcd_clk,
    kcd_reset       => kcd_reset,
    cmd_valid       => sum_base_price_inst_cmd_valid,
    cmd_ready       => sum_base_price_inst_cmd_ready,
    cmd_firstIdx    => sum_base_price_inst_cmd_firstIdx,
    cmd_lastIdx     => sum_base_price_inst_cmd_lastIdx,
    cmd_ctrl        => sum_base_price_inst_cmd_ctrl,
    cmd_tag         => sum_base_price_inst_cmd_tag,
    unl_valid       => sum_base_price_inst_unl_valid,
    unl_ready       => sum_base_price_inst_unl_ready,
    unl_tag         => sum_base_price_inst_unl_tag,
    bus_wreq_valid  => sum_base_price_inst_bus_wreq_valid,
    bus_wreq_ready  => sum_base_price_inst_bus_wreq_ready,
    bus_wreq_addr   => sum_base_price_inst_bus_wreq_addr,
    bus_wreq_len    => sum_base_price_inst_bus_wreq_len,
    bus_wreq_last   => sum_base_price_inst_bus_wreq_last,
    bus_wdat_valid  => sum_base_price_inst_bus_wdat_valid,
    bus_wdat_ready  => sum_base_price_inst_bus_wdat_ready,
    bus_wdat_data   => sum_base_price_inst_bus_wdat_data,
    bus_wdat_strobe => sum_base_price_inst_bus_wdat_strobe,
    bus_wdat_last   => sum_base_price_inst_bus_wdat_last,
    bus_wrep_valid  => sum_base_price_inst_bus_wrep_valid,
    bus_wrep_ready  => sum_base_price_inst_bus_wrep_ready,
    bus_wrep_ok     => sum_base_price_inst_bus_wrep_ok,
    in_valid        => sum_base_price_inst_in_valid,
    in_ready        => sum_base_price_inst_in_ready,
    in_data         => sum_base_price_inst_in_data,
    in_dvalid       => sum_base_price_inst_in_dvalid,
    in_last         => sum_base_price_inst_in_last
  );

  sum_disc_price_inst : ArrayWriter
  generic map(
    BUS_ADDR_WIDTH     => L_SUM_DISC_PRICE_BUS_ADDR_WIDTH,
    BUS_DATA_WIDTH     => L_SUM_DISC_PRICE_BUS_DATA_WIDTH,
    BUS_LEN_WIDTH      => L_SUM_DISC_PRICE_BUS_LEN_WIDTH,
    BUS_BURST_STEP_LEN => L_SUM_DISC_PRICE_BUS_BURST_STEP_LEN,
    BUS_BURST_MAX_LEN  => L_SUM_DISC_PRICE_BUS_BURST_MAX_LEN,
    INDEX_WIDTH        => INDEX_WIDTH,
    CFG                => "prim(64)",
    CMD_TAG_ENABLE     => true,
    CMD_TAG_WIDTH      => TAG_WIDTH
  )
  port map(
    bcd_clk         => bcd_clk,
    bcd_reset       => bcd_reset,
    kcd_clk         => kcd_clk,
    kcd_reset       => kcd_reset,
    cmd_valid       => sum_disc_price_inst_cmd_valid,
    cmd_ready       => sum_disc_price_inst_cmd_ready,
    cmd_firstIdx    => sum_disc_price_inst_cmd_firstIdx,
    cmd_lastIdx     => sum_disc_price_inst_cmd_lastIdx,
    cmd_ctrl        => sum_disc_price_inst_cmd_ctrl,
    cmd_tag         => sum_disc_price_inst_cmd_tag,
    unl_valid       => sum_disc_price_inst_unl_valid,
    unl_ready       => sum_disc_price_inst_unl_ready,
    unl_tag         => sum_disc_price_inst_unl_tag,
    bus_wreq_valid  => sum_disc_price_inst_bus_wreq_valid,
    bus_wreq_ready  => sum_disc_price_inst_bus_wreq_ready,
    bus_wreq_addr   => sum_disc_price_inst_bus_wreq_addr,
    bus_wreq_len    => sum_disc_price_inst_bus_wreq_len,
    bus_wreq_last   => sum_disc_price_inst_bus_wreq_last,
    bus_wdat_valid  => sum_disc_price_inst_bus_wdat_valid,
    bus_wdat_ready  => sum_disc_price_inst_bus_wdat_ready,
    bus_wdat_data   => sum_disc_price_inst_bus_wdat_data,
    bus_wdat_strobe => sum_disc_price_inst_bus_wdat_strobe,
    bus_wdat_last   => sum_disc_price_inst_bus_wdat_last,
    bus_wrep_valid  => sum_disc_price_inst_bus_wrep_valid,
    bus_wrep_ready  => sum_disc_price_inst_bus_wrep_ready,
    bus_wrep_ok     => sum_disc_price_inst_bus_wrep_ok,
    in_valid        => sum_disc_price_inst_in_valid,
    in_ready        => sum_disc_price_inst_in_ready,
    in_data         => sum_disc_price_inst_in_data,
    in_dvalid       => sum_disc_price_inst_in_dvalid,
    in_last         => sum_disc_price_inst_in_last
  );

  sum_charge_inst : ArrayWriter
  generic map(
    BUS_ADDR_WIDTH     => L_SUM_CHARGE_BUS_ADDR_WIDTH,
    BUS_DATA_WIDTH     => L_SUM_CHARGE_BUS_DATA_WIDTH,
    BUS_LEN_WIDTH      => L_SUM_CHARGE_BUS_LEN_WIDTH,
    BUS_BURST_STEP_LEN => L_SUM_CHARGE_BUS_BURST_STEP_LEN,
    BUS_BURST_MAX_LEN  => L_SUM_CHARGE_BUS_BURST_MAX_LEN,
    INDEX_WIDTH        => INDEX_WIDTH,
    CFG                => "prim(64)",
    CMD_TAG_ENABLE     => true,
    CMD_TAG_WIDTH      => TAG_WIDTH
  )
  port map(
    bcd_clk         => bcd_clk,
    bcd_reset       => bcd_reset,
    kcd_clk         => kcd_clk,
    kcd_reset       => kcd_reset,
    cmd_valid       => sum_charge_inst_cmd_valid,
    cmd_ready       => sum_charge_inst_cmd_ready,
    cmd_firstIdx    => sum_charge_inst_cmd_firstIdx,
    cmd_lastIdx     => sum_charge_inst_cmd_lastIdx,
    cmd_ctrl        => sum_charge_inst_cmd_ctrl,
    cmd_tag         => sum_charge_inst_cmd_tag,
    unl_valid       => sum_charge_inst_unl_valid,
    unl_ready       => sum_charge_inst_unl_ready,
    unl_tag         => sum_charge_inst_unl_tag,
    bus_wreq_valid  => sum_charge_inst_bus_wreq_valid,
    bus_wreq_ready  => sum_charge_inst_bus_wreq_ready,
    bus_wreq_addr   => sum_charge_inst_bus_wreq_addr,
    bus_wreq_len    => sum_charge_inst_bus_wreq_len,
    bus_wreq_last   => sum_charge_inst_bus_wreq_last,
    bus_wdat_valid  => sum_charge_inst_bus_wdat_valid,
    bus_wdat_ready  => sum_charge_inst_bus_wdat_ready,
    bus_wdat_data   => sum_charge_inst_bus_wdat_data,
    bus_wdat_strobe => sum_charge_inst_bus_wdat_strobe,
    bus_wdat_last   => sum_charge_inst_bus_wdat_last,
    bus_wrep_valid  => sum_charge_inst_bus_wrep_valid,
    bus_wrep_ready  => sum_charge_inst_bus_wrep_ready,
    bus_wrep_ok     => sum_charge_inst_bus_wrep_ok,
    in_valid        => sum_charge_inst_in_valid,
    in_ready        => sum_charge_inst_in_ready,
    in_data         => sum_charge_inst_in_data,
    in_dvalid       => sum_charge_inst_in_dvalid,
    in_last         => sum_charge_inst_in_last
  );

  avg_qty_inst : ArrayWriter
  generic map(
    BUS_ADDR_WIDTH     => L_AVG_QTY_BUS_ADDR_WIDTH,
    BUS_DATA_WIDTH     => L_AVG_QTY_BUS_DATA_WIDTH,
    BUS_LEN_WIDTH      => L_AVG_QTY_BUS_LEN_WIDTH,
    BUS_BURST_STEP_LEN => L_AVG_QTY_BUS_BURST_STEP_LEN,
    BUS_BURST_MAX_LEN  => L_AVG_QTY_BUS_BURST_MAX_LEN,
    INDEX_WIDTH        => INDEX_WIDTH,
    CFG                => "prim(64)",
    CMD_TAG_ENABLE     => true,
    CMD_TAG_WIDTH      => TAG_WIDTH
  )
  port map(
    bcd_clk         => bcd_clk,
    bcd_reset       => bcd_reset,
    kcd_clk         => kcd_clk,
    kcd_reset       => kcd_reset,
    cmd_valid       => avg_qty_inst_cmd_valid,
    cmd_ready       => avg_qty_inst_cmd_ready,
    cmd_firstIdx    => avg_qty_inst_cmd_firstIdx,
    cmd_lastIdx     => avg_qty_inst_cmd_lastIdx,
    cmd_ctrl        => avg_qty_inst_cmd_ctrl,
    cmd_tag         => avg_qty_inst_cmd_tag,
    unl_valid       => avg_qty_inst_unl_valid,
    unl_ready       => avg_qty_inst_unl_ready,
    unl_tag         => avg_qty_inst_unl_tag,
    bus_wreq_valid  => avg_qty_inst_bus_wreq_valid,
    bus_wreq_ready  => avg_qty_inst_bus_wreq_ready,
    bus_wreq_addr   => avg_qty_inst_bus_wreq_addr,
    bus_wreq_len    => avg_qty_inst_bus_wreq_len,
    bus_wreq_last   => avg_qty_inst_bus_wreq_last,
    bus_wdat_valid  => avg_qty_inst_bus_wdat_valid,
    bus_wdat_ready  => avg_qty_inst_bus_wdat_ready,
    bus_wdat_data   => avg_qty_inst_bus_wdat_data,
    bus_wdat_strobe => avg_qty_inst_bus_wdat_strobe,
    bus_wdat_last   => avg_qty_inst_bus_wdat_last,
    bus_wrep_valid  => avg_qty_inst_bus_wrep_valid,
    bus_wrep_ready  => avg_qty_inst_bus_wrep_ready,
    bus_wrep_ok     => avg_qty_inst_bus_wrep_ok,
    in_valid        => avg_qty_inst_in_valid,
    in_ready        => avg_qty_inst_in_ready,
    in_data         => avg_qty_inst_in_data,
    in_dvalid       => avg_qty_inst_in_dvalid,
    in_last         => avg_qty_inst_in_last
  );

  avg_price_inst : ArrayWriter
  generic map(
    BUS_ADDR_WIDTH     => L_AVG_PRICE_BUS_ADDR_WIDTH,
    BUS_DATA_WIDTH     => L_AVG_PRICE_BUS_DATA_WIDTH,
    BUS_LEN_WIDTH      => L_AVG_PRICE_BUS_LEN_WIDTH,
    BUS_BURST_STEP_LEN => L_AVG_PRICE_BUS_BURST_STEP_LEN,
    BUS_BURST_MAX_LEN  => L_AVG_PRICE_BUS_BURST_MAX_LEN,
    INDEX_WIDTH        => INDEX_WIDTH,
    CFG                => "prim(64)",
    CMD_TAG_ENABLE     => true,
    CMD_TAG_WIDTH      => TAG_WIDTH
  )
  port map(
    bcd_clk         => bcd_clk,
    bcd_reset       => bcd_reset,
    kcd_clk         => kcd_clk,
    kcd_reset       => kcd_reset,
    cmd_valid       => avg_price_inst_cmd_valid,
    cmd_ready       => avg_price_inst_cmd_ready,
    cmd_firstIdx    => avg_price_inst_cmd_firstIdx,
    cmd_lastIdx     => avg_price_inst_cmd_lastIdx,
    cmd_ctrl        => avg_price_inst_cmd_ctrl,
    cmd_tag         => avg_price_inst_cmd_tag,
    unl_valid       => avg_price_inst_unl_valid,
    unl_ready       => avg_price_inst_unl_ready,
    unl_tag         => avg_price_inst_unl_tag,
    bus_wreq_valid  => avg_price_inst_bus_wreq_valid,
    bus_wreq_ready  => avg_price_inst_bus_wreq_ready,
    bus_wreq_addr   => avg_price_inst_bus_wreq_addr,
    bus_wreq_len    => avg_price_inst_bus_wreq_len,
    bus_wreq_last   => avg_price_inst_bus_wreq_last,
    bus_wdat_valid  => avg_price_inst_bus_wdat_valid,
    bus_wdat_ready  => avg_price_inst_bus_wdat_ready,
    bus_wdat_data   => avg_price_inst_bus_wdat_data,
    bus_wdat_strobe => avg_price_inst_bus_wdat_strobe,
    bus_wdat_last   => avg_price_inst_bus_wdat_last,
    bus_wrep_valid  => avg_price_inst_bus_wrep_valid,
    bus_wrep_ready  => avg_price_inst_bus_wrep_ready,
    bus_wrep_ok     => avg_price_inst_bus_wrep_ok,
    in_valid        => avg_price_inst_in_valid,
    in_ready        => avg_price_inst_in_ready,
    in_data         => avg_price_inst_in_data,
    in_dvalid       => avg_price_inst_in_dvalid,
    in_last         => avg_price_inst_in_last
  );

  avg_disc_inst : ArrayWriter
  generic map(
    BUS_ADDR_WIDTH     => L_AVG_DISC_BUS_ADDR_WIDTH,
    BUS_DATA_WIDTH     => L_AVG_DISC_BUS_DATA_WIDTH,
    BUS_LEN_WIDTH      => L_AVG_DISC_BUS_LEN_WIDTH,
    BUS_BURST_STEP_LEN => L_AVG_DISC_BUS_BURST_STEP_LEN,
    BUS_BURST_MAX_LEN  => L_AVG_DISC_BUS_BURST_MAX_LEN,
    INDEX_WIDTH        => INDEX_WIDTH,
    CFG                => "prim(64)",
    CMD_TAG_ENABLE     => true,
    CMD_TAG_WIDTH      => TAG_WIDTH
  )
  port map(
    bcd_clk         => bcd_clk,
    bcd_reset       => bcd_reset,
    kcd_clk         => kcd_clk,
    kcd_reset       => kcd_reset,
    cmd_valid       => avg_disc_inst_cmd_valid,
    cmd_ready       => avg_disc_inst_cmd_ready,
    cmd_firstIdx    => avg_disc_inst_cmd_firstIdx,
    cmd_lastIdx     => avg_disc_inst_cmd_lastIdx,
    cmd_ctrl        => avg_disc_inst_cmd_ctrl,
    cmd_tag         => avg_disc_inst_cmd_tag,
    unl_valid       => avg_disc_inst_unl_valid,
    unl_ready       => avg_disc_inst_unl_ready,
    unl_tag         => avg_disc_inst_unl_tag,
    bus_wreq_valid  => avg_disc_inst_bus_wreq_valid,
    bus_wreq_ready  => avg_disc_inst_bus_wreq_ready,
    bus_wreq_addr   => avg_disc_inst_bus_wreq_addr,
    bus_wreq_len    => avg_disc_inst_bus_wreq_len,
    bus_wreq_last   => avg_disc_inst_bus_wreq_last,
    bus_wdat_valid  => avg_disc_inst_bus_wdat_valid,
    bus_wdat_ready  => avg_disc_inst_bus_wdat_ready,
    bus_wdat_data   => avg_disc_inst_bus_wdat_data,
    bus_wdat_strobe => avg_disc_inst_bus_wdat_strobe,
    bus_wdat_last   => avg_disc_inst_bus_wdat_last,
    bus_wrep_valid  => avg_disc_inst_bus_wrep_valid,
    bus_wrep_ready  => avg_disc_inst_bus_wrep_ready,
    bus_wrep_ok     => avg_disc_inst_bus_wrep_ok,
    in_valid        => avg_disc_inst_in_valid,
    in_ready        => avg_disc_inst_in_ready,
    in_data         => avg_disc_inst_in_data,
    in_dvalid       => avg_disc_inst_in_dvalid,
    in_last         => avg_disc_inst_in_last
  );

  count_order_inst : ArrayWriter
  generic map(
    BUS_ADDR_WIDTH     => L_COUNT_ORDER_BUS_ADDR_WIDTH,
    BUS_DATA_WIDTH     => L_COUNT_ORDER_BUS_DATA_WIDTH,
    BUS_LEN_WIDTH      => L_COUNT_ORDER_BUS_LEN_WIDTH,
    BUS_BURST_STEP_LEN => L_COUNT_ORDER_BUS_BURST_STEP_LEN,
    BUS_BURST_MAX_LEN  => L_COUNT_ORDER_BUS_BURST_MAX_LEN,
    INDEX_WIDTH        => INDEX_WIDTH,
    CFG                => "prim(64)",
    CMD_TAG_ENABLE     => true,
    CMD_TAG_WIDTH      => TAG_WIDTH
  )
  port map(
    bcd_clk         => bcd_clk,
    bcd_reset       => bcd_reset,
    kcd_clk         => kcd_clk,
    kcd_reset       => kcd_reset,
    cmd_valid       => count_order_inst_cmd_valid,
    cmd_ready       => count_order_inst_cmd_ready,
    cmd_firstIdx    => count_order_inst_cmd_firstIdx,
    cmd_lastIdx     => count_order_inst_cmd_lastIdx,
    cmd_ctrl        => count_order_inst_cmd_ctrl,
    cmd_tag         => count_order_inst_cmd_tag,
    unl_valid       => count_order_inst_unl_valid,
    unl_ready       => count_order_inst_unl_ready,
    unl_tag         => count_order_inst_unl_tag,
    bus_wreq_valid  => count_order_inst_bus_wreq_valid,
    bus_wreq_ready  => count_order_inst_bus_wreq_ready,
    bus_wreq_addr   => count_order_inst_bus_wreq_addr,
    bus_wreq_len    => count_order_inst_bus_wreq_len,
    bus_wreq_last   => count_order_inst_bus_wreq_last,
    bus_wdat_valid  => count_order_inst_bus_wdat_valid,
    bus_wdat_ready  => count_order_inst_bus_wdat_ready,
    bus_wdat_data   => count_order_inst_bus_wdat_data,
    bus_wdat_strobe => count_order_inst_bus_wdat_strobe,
    bus_wdat_last   => count_order_inst_bus_wdat_last,
    bus_wrep_valid  => count_order_inst_bus_wrep_valid,
    bus_wrep_ready  => count_order_inst_bus_wrep_ready,
    bus_wrep_ok     => count_order_inst_bus_wrep_ok,
    in_valid        => count_order_inst_in_valid,
    in_ready        => count_order_inst_in_ready,
    in_data         => count_order_inst_in_data,
    in_dvalid       => count_order_inst_in_dvalid,
    in_last         => count_order_inst_in_last
  );

  l_returnflag_o_bus_wreq_valid           <= returnflag_o_inst_bus_wreq_valid;
  returnflag_o_inst_bus_wreq_ready        <= l_returnflag_o_bus_wreq_ready;
  l_returnflag_o_bus_wreq_addr            <= returnflag_o_inst_bus_wreq_addr;
  l_returnflag_o_bus_wreq_len             <= returnflag_o_inst_bus_wreq_len;
  l_returnflag_o_bus_wreq_last            <= returnflag_o_inst_bus_wreq_last;
  l_returnflag_o_bus_wdat_valid           <= returnflag_o_inst_bus_wdat_valid;
  returnflag_o_inst_bus_wdat_ready        <= l_returnflag_o_bus_wdat_ready;
  l_returnflag_o_bus_wdat_data            <= returnflag_o_inst_bus_wdat_data;
  l_returnflag_o_bus_wdat_strobe          <= returnflag_o_inst_bus_wdat_strobe;
  l_returnflag_o_bus_wdat_last            <= returnflag_o_inst_bus_wdat_last;
  returnflag_o_inst_bus_wrep_valid        <= l_returnflag_o_bus_wrep_valid;
  l_returnflag_o_bus_wrep_ready           <= returnflag_o_inst_bus_wrep_ready;
  returnflag_o_inst_bus_wrep_ok           <= l_returnflag_o_bus_wrep_ok;

  l_returnflag_o_unl_valid                <= returnflag_o_inst_unl_valid;
  returnflag_o_inst_unl_ready             <= l_returnflag_o_unl_ready;
  l_returnflag_o_unl_tag                  <= returnflag_o_inst_unl_tag;

  l_linestatus_o_bus_wreq_valid           <= linestatus_o_inst_bus_wreq_valid;
  linestatus_o_inst_bus_wreq_ready        <= l_linestatus_o_bus_wreq_ready;
  l_linestatus_o_bus_wreq_addr            <= linestatus_o_inst_bus_wreq_addr;
  l_linestatus_o_bus_wreq_len             <= linestatus_o_inst_bus_wreq_len;
  l_linestatus_o_bus_wreq_last            <= linestatus_o_inst_bus_wreq_last;
  l_linestatus_o_bus_wdat_valid           <= linestatus_o_inst_bus_wdat_valid;
  linestatus_o_inst_bus_wdat_ready        <= l_linestatus_o_bus_wdat_ready;
  l_linestatus_o_bus_wdat_data            <= linestatus_o_inst_bus_wdat_data;
  l_linestatus_o_bus_wdat_strobe          <= linestatus_o_inst_bus_wdat_strobe;
  l_linestatus_o_bus_wdat_last            <= linestatus_o_inst_bus_wdat_last;
  linestatus_o_inst_bus_wrep_valid        <= l_linestatus_o_bus_wrep_valid;
  l_linestatus_o_bus_wrep_ready           <= linestatus_o_inst_bus_wrep_ready;
  linestatus_o_inst_bus_wrep_ok           <= l_linestatus_o_bus_wrep_ok;

  l_linestatus_o_unl_valid                <= linestatus_o_inst_unl_valid;
  linestatus_o_inst_unl_ready             <= l_linestatus_o_unl_ready;
  l_linestatus_o_unl_tag                  <= linestatus_o_inst_unl_tag;

  l_sum_qty_bus_wreq_valid                <= sum_qty_inst_bus_wreq_valid;
  sum_qty_inst_bus_wreq_ready             <= l_sum_qty_bus_wreq_ready;
  l_sum_qty_bus_wreq_addr                 <= sum_qty_inst_bus_wreq_addr;
  l_sum_qty_bus_wreq_len                  <= sum_qty_inst_bus_wreq_len;
  l_sum_qty_bus_wreq_last                 <= sum_qty_inst_bus_wreq_last;
  l_sum_qty_bus_wdat_valid                <= sum_qty_inst_bus_wdat_valid;
  sum_qty_inst_bus_wdat_ready             <= l_sum_qty_bus_wdat_ready;
  l_sum_qty_bus_wdat_data                 <= sum_qty_inst_bus_wdat_data;
  l_sum_qty_bus_wdat_strobe               <= sum_qty_inst_bus_wdat_strobe;
  l_sum_qty_bus_wdat_last                 <= sum_qty_inst_bus_wdat_last;
  sum_qty_inst_bus_wrep_valid             <= l_sum_qty_bus_wrep_valid;
  l_sum_qty_bus_wrep_ready                <= sum_qty_inst_bus_wrep_ready;
  sum_qty_inst_bus_wrep_ok                <= l_sum_qty_bus_wrep_ok;

  l_sum_qty_unl_valid                     <= sum_qty_inst_unl_valid;
  sum_qty_inst_unl_ready                  <= l_sum_qty_unl_ready;
  l_sum_qty_unl_tag                       <= sum_qty_inst_unl_tag;

  l_sum_base_price_bus_wreq_valid         <= sum_base_price_inst_bus_wreq_valid;
  sum_base_price_inst_bus_wreq_ready      <= l_sum_base_price_bus_wreq_ready;
  l_sum_base_price_bus_wreq_addr          <= sum_base_price_inst_bus_wreq_addr;
  l_sum_base_price_bus_wreq_len           <= sum_base_price_inst_bus_wreq_len;
  l_sum_base_price_bus_wreq_last          <= sum_base_price_inst_bus_wreq_last;
  l_sum_base_price_bus_wdat_valid         <= sum_base_price_inst_bus_wdat_valid;
  sum_base_price_inst_bus_wdat_ready      <= l_sum_base_price_bus_wdat_ready;
  l_sum_base_price_bus_wdat_data          <= sum_base_price_inst_bus_wdat_data;
  l_sum_base_price_bus_wdat_strobe        <= sum_base_price_inst_bus_wdat_strobe;
  l_sum_base_price_bus_wdat_last          <= sum_base_price_inst_bus_wdat_last;
  sum_base_price_inst_bus_wrep_valid      <= l_sum_base_price_bus_wrep_valid;
  l_sum_base_price_bus_wrep_ready         <= sum_base_price_inst_bus_wrep_ready;
  sum_base_price_inst_bus_wrep_ok         <= l_sum_base_price_bus_wrep_ok;

  l_sum_base_price_unl_valid              <= sum_base_price_inst_unl_valid;
  sum_base_price_inst_unl_ready           <= l_sum_base_price_unl_ready;
  l_sum_base_price_unl_tag                <= sum_base_price_inst_unl_tag;

  l_sum_disc_price_bus_wreq_valid         <= sum_disc_price_inst_bus_wreq_valid;
  sum_disc_price_inst_bus_wreq_ready      <= l_sum_disc_price_bus_wreq_ready;
  l_sum_disc_price_bus_wreq_addr          <= sum_disc_price_inst_bus_wreq_addr;
  l_sum_disc_price_bus_wreq_len           <= sum_disc_price_inst_bus_wreq_len;
  l_sum_disc_price_bus_wreq_last          <= sum_disc_price_inst_bus_wreq_last;
  l_sum_disc_price_bus_wdat_valid         <= sum_disc_price_inst_bus_wdat_valid;
  sum_disc_price_inst_bus_wdat_ready      <= l_sum_disc_price_bus_wdat_ready;
  l_sum_disc_price_bus_wdat_data          <= sum_disc_price_inst_bus_wdat_data;
  l_sum_disc_price_bus_wdat_strobe        <= sum_disc_price_inst_bus_wdat_strobe;
  l_sum_disc_price_bus_wdat_last          <= sum_disc_price_inst_bus_wdat_last;
  sum_disc_price_inst_bus_wrep_valid      <= l_sum_disc_price_bus_wrep_valid;
  l_sum_disc_price_bus_wrep_ready         <= sum_disc_price_inst_bus_wrep_ready;
  sum_disc_price_inst_bus_wrep_ok         <= l_sum_disc_price_bus_wrep_ok;

  l_sum_disc_price_unl_valid              <= sum_disc_price_inst_unl_valid;
  sum_disc_price_inst_unl_ready           <= l_sum_disc_price_unl_ready;
  l_sum_disc_price_unl_tag                <= sum_disc_price_inst_unl_tag;

  l_sum_charge_bus_wreq_valid             <= sum_charge_inst_bus_wreq_valid;
  sum_charge_inst_bus_wreq_ready          <= l_sum_charge_bus_wreq_ready;
  l_sum_charge_bus_wreq_addr              <= sum_charge_inst_bus_wreq_addr;
  l_sum_charge_bus_wreq_len               <= sum_charge_inst_bus_wreq_len;
  l_sum_charge_bus_wreq_last              <= sum_charge_inst_bus_wreq_last;
  l_sum_charge_bus_wdat_valid             <= sum_charge_inst_bus_wdat_valid;
  sum_charge_inst_bus_wdat_ready          <= l_sum_charge_bus_wdat_ready;
  l_sum_charge_bus_wdat_data              <= sum_charge_inst_bus_wdat_data;
  l_sum_charge_bus_wdat_strobe            <= sum_charge_inst_bus_wdat_strobe;
  l_sum_charge_bus_wdat_last              <= sum_charge_inst_bus_wdat_last;
  sum_charge_inst_bus_wrep_valid          <= l_sum_charge_bus_wrep_valid;
  l_sum_charge_bus_wrep_ready             <= sum_charge_inst_bus_wrep_ready;
  sum_charge_inst_bus_wrep_ok             <= l_sum_charge_bus_wrep_ok;

  l_sum_charge_unl_valid                  <= sum_charge_inst_unl_valid;
  sum_charge_inst_unl_ready               <= l_sum_charge_unl_ready;
  l_sum_charge_unl_tag                    <= sum_charge_inst_unl_tag;

  l_avg_qty_bus_wreq_valid                <= avg_qty_inst_bus_wreq_valid;
  avg_qty_inst_bus_wreq_ready             <= l_avg_qty_bus_wreq_ready;
  l_avg_qty_bus_wreq_addr                 <= avg_qty_inst_bus_wreq_addr;
  l_avg_qty_bus_wreq_len                  <= avg_qty_inst_bus_wreq_len;
  l_avg_qty_bus_wreq_last                 <= avg_qty_inst_bus_wreq_last;
  l_avg_qty_bus_wdat_valid                <= avg_qty_inst_bus_wdat_valid;
  avg_qty_inst_bus_wdat_ready             <= l_avg_qty_bus_wdat_ready;
  l_avg_qty_bus_wdat_data                 <= avg_qty_inst_bus_wdat_data;
  l_avg_qty_bus_wdat_strobe               <= avg_qty_inst_bus_wdat_strobe;
  l_avg_qty_bus_wdat_last                 <= avg_qty_inst_bus_wdat_last;
  avg_qty_inst_bus_wrep_valid             <= l_avg_qty_bus_wrep_valid;
  l_avg_qty_bus_wrep_ready                <= avg_qty_inst_bus_wrep_ready;
  avg_qty_inst_bus_wrep_ok                <= l_avg_qty_bus_wrep_ok;

  l_avg_qty_unl_valid                     <= avg_qty_inst_unl_valid;
  avg_qty_inst_unl_ready                  <= l_avg_qty_unl_ready;
  l_avg_qty_unl_tag                       <= avg_qty_inst_unl_tag;

  l_avg_price_bus_wreq_valid              <= avg_price_inst_bus_wreq_valid;
  avg_price_inst_bus_wreq_ready           <= l_avg_price_bus_wreq_ready;
  l_avg_price_bus_wreq_addr               <= avg_price_inst_bus_wreq_addr;
  l_avg_price_bus_wreq_len                <= avg_price_inst_bus_wreq_len;
  l_avg_price_bus_wreq_last               <= avg_price_inst_bus_wreq_last;
  l_avg_price_bus_wdat_valid              <= avg_price_inst_bus_wdat_valid;
  avg_price_inst_bus_wdat_ready           <= l_avg_price_bus_wdat_ready;
  l_avg_price_bus_wdat_data               <= avg_price_inst_bus_wdat_data;
  l_avg_price_bus_wdat_strobe             <= avg_price_inst_bus_wdat_strobe;
  l_avg_price_bus_wdat_last               <= avg_price_inst_bus_wdat_last;
  avg_price_inst_bus_wrep_valid           <= l_avg_price_bus_wrep_valid;
  l_avg_price_bus_wrep_ready              <= avg_price_inst_bus_wrep_ready;
  avg_price_inst_bus_wrep_ok              <= l_avg_price_bus_wrep_ok;

  l_avg_price_unl_valid                   <= avg_price_inst_unl_valid;
  avg_price_inst_unl_ready                <= l_avg_price_unl_ready;
  l_avg_price_unl_tag                     <= avg_price_inst_unl_tag;

  l_avg_disc_bus_wreq_valid               <= avg_disc_inst_bus_wreq_valid;
  avg_disc_inst_bus_wreq_ready            <= l_avg_disc_bus_wreq_ready;
  l_avg_disc_bus_wreq_addr                <= avg_disc_inst_bus_wreq_addr;
  l_avg_disc_bus_wreq_len                 <= avg_disc_inst_bus_wreq_len;
  l_avg_disc_bus_wreq_last                <= avg_disc_inst_bus_wreq_last;
  l_avg_disc_bus_wdat_valid               <= avg_disc_inst_bus_wdat_valid;
  avg_disc_inst_bus_wdat_ready            <= l_avg_disc_bus_wdat_ready;
  l_avg_disc_bus_wdat_data                <= avg_disc_inst_bus_wdat_data;
  l_avg_disc_bus_wdat_strobe              <= avg_disc_inst_bus_wdat_strobe;
  l_avg_disc_bus_wdat_last                <= avg_disc_inst_bus_wdat_last;
  avg_disc_inst_bus_wrep_valid            <= l_avg_disc_bus_wrep_valid;
  l_avg_disc_bus_wrep_ready               <= avg_disc_inst_bus_wrep_ready;
  avg_disc_inst_bus_wrep_ok               <= l_avg_disc_bus_wrep_ok;

  l_avg_disc_unl_valid                    <= avg_disc_inst_unl_valid;
  avg_disc_inst_unl_ready                 <= l_avg_disc_unl_ready;
  l_avg_disc_unl_tag                      <= avg_disc_inst_unl_tag;

  l_count_order_bus_wreq_valid            <= count_order_inst_bus_wreq_valid;
  count_order_inst_bus_wreq_ready         <= l_count_order_bus_wreq_ready;
  l_count_order_bus_wreq_addr             <= count_order_inst_bus_wreq_addr;
  l_count_order_bus_wreq_len              <= count_order_inst_bus_wreq_len;
  l_count_order_bus_wreq_last             <= count_order_inst_bus_wreq_last;
  l_count_order_bus_wdat_valid            <= count_order_inst_bus_wdat_valid;
  count_order_inst_bus_wdat_ready         <= l_count_order_bus_wdat_ready;
  l_count_order_bus_wdat_data             <= count_order_inst_bus_wdat_data;
  l_count_order_bus_wdat_strobe           <= count_order_inst_bus_wdat_strobe;
  l_count_order_bus_wdat_last             <= count_order_inst_bus_wdat_last;
  count_order_inst_bus_wrep_valid         <= l_count_order_bus_wrep_valid;
  l_count_order_bus_wrep_ready            <= count_order_inst_bus_wrep_ready;
  count_order_inst_bus_wrep_ok            <= l_count_order_bus_wrep_ok;

  l_count_order_unl_valid                 <= count_order_inst_unl_valid;
  count_order_inst_unl_ready              <= l_count_order_unl_ready;
  l_count_order_unl_tag                   <= count_order_inst_unl_tag;

  returnflag_o_inst_cmd_valid             <= l_returnflag_o_cmd_valid;
  l_returnflag_o_cmd_ready                <= returnflag_o_inst_cmd_ready;
  returnflag_o_inst_cmd_firstIdx          <= l_returnflag_o_cmd_firstIdx;
  returnflag_o_inst_cmd_lastIdx           <= l_returnflag_o_cmd_lastIdx;
  returnflag_o_inst_cmd_ctrl              <= l_returnflag_o_cmd_ctrl;
  returnflag_o_inst_cmd_tag               <= l_returnflag_o_cmd_tag;

  returnflag_o_inst_in_valid(0)           <= l_returnflag_o_valid;
  returnflag_o_inst_in_valid(1)           <= l_returnflag_o_chars_valid;
  l_returnflag_o_ready                    <= returnflag_o_inst_in_ready(0);
  l_returnflag_o_chars_ready              <= returnflag_o_inst_in_ready(1);
  returnflag_o_inst_in_data(31 downto 0)  <= l_returnflag_o_length;
  returnflag_o_inst_in_data(32 downto 32) <= l_returnflag_o_count;
  returnflag_o_inst_in_data(40 downto 33) <= l_returnflag_o_chars;
  returnflag_o_inst_in_data(41 downto 41) <= l_returnflag_o_chars_count;
  returnflag_o_inst_in_dvalid(0)          <= l_returnflag_o_dvalid;
  returnflag_o_inst_in_dvalid(1)          <= l_returnflag_o_chars_dvalid;
  returnflag_o_inst_in_last(0)            <= l_returnflag_o_last;
  returnflag_o_inst_in_last(1)            <= l_returnflag_o_chars_last;

  linestatus_o_inst_cmd_valid             <= l_linestatus_o_cmd_valid;
  l_linestatus_o_cmd_ready                <= linestatus_o_inst_cmd_ready;
  linestatus_o_inst_cmd_firstIdx          <= l_linestatus_o_cmd_firstIdx;
  linestatus_o_inst_cmd_lastIdx           <= l_linestatus_o_cmd_lastIdx;
  linestatus_o_inst_cmd_ctrl              <= l_linestatus_o_cmd_ctrl;
  linestatus_o_inst_cmd_tag               <= l_linestatus_o_cmd_tag;

  linestatus_o_inst_in_valid(0)           <= l_linestatus_o_valid;
  linestatus_o_inst_in_valid(1)           <= l_linestatus_o_chars_valid;
  l_linestatus_o_ready                    <= linestatus_o_inst_in_ready(0);
  l_linestatus_o_chars_ready              <= linestatus_o_inst_in_ready(1);
  linestatus_o_inst_in_data(31 downto 0)  <= l_linestatus_o_length;
  linestatus_o_inst_in_data(32 downto 32) <= l_linestatus_o_count;
  linestatus_o_inst_in_data(40 downto 33) <= l_linestatus_o_chars;
  linestatus_o_inst_in_data(41 downto 41) <= l_linestatus_o_chars_count;
  linestatus_o_inst_in_dvalid(0)          <= l_linestatus_o_dvalid;
  linestatus_o_inst_in_dvalid(1)          <= l_linestatus_o_chars_dvalid;
  linestatus_o_inst_in_last(0)            <= l_linestatus_o_last;
  linestatus_o_inst_in_last(1)            <= l_linestatus_o_chars_last;

  sum_qty_inst_cmd_valid                  <= l_sum_qty_cmd_valid;
  l_sum_qty_cmd_ready                     <= sum_qty_inst_cmd_ready;
  sum_qty_inst_cmd_firstIdx               <= l_sum_qty_cmd_firstIdx;
  sum_qty_inst_cmd_lastIdx                <= l_sum_qty_cmd_lastIdx;
  sum_qty_inst_cmd_ctrl                   <= l_sum_qty_cmd_ctrl;
  sum_qty_inst_cmd_tag                    <= l_sum_qty_cmd_tag;

  sum_qty_inst_in_valid(0)                <= l_sum_qty_valid;
  l_sum_qty_ready                         <= sum_qty_inst_in_ready(0);
  sum_qty_inst_in_data                    <= l_sum_qty;
  sum_qty_inst_in_dvalid(0)               <= l_sum_qty_dvalid;
  sum_qty_inst_in_last(0)                 <= l_sum_qty_last;

  sum_base_price_inst_cmd_valid           <= l_sum_base_price_cmd_valid;
  l_sum_base_price_cmd_ready              <= sum_base_price_inst_cmd_ready;
  sum_base_price_inst_cmd_firstIdx        <= l_sum_base_price_cmd_firstIdx;
  sum_base_price_inst_cmd_lastIdx         <= l_sum_base_price_cmd_lastIdx;
  sum_base_price_inst_cmd_ctrl            <= l_sum_base_price_cmd_ctrl;
  sum_base_price_inst_cmd_tag             <= l_sum_base_price_cmd_tag;

  sum_base_price_inst_in_valid(0)         <= l_sum_base_price_valid;
  l_sum_base_price_ready                  <= sum_base_price_inst_in_ready(0);
  sum_base_price_inst_in_data             <= l_sum_base_price;
  sum_base_price_inst_in_dvalid(0)        <= l_sum_base_price_dvalid;
  sum_base_price_inst_in_last(0)          <= l_sum_base_price_last;

  sum_disc_price_inst_cmd_valid           <= l_sum_disc_price_cmd_valid;
  l_sum_disc_price_cmd_ready              <= sum_disc_price_inst_cmd_ready;
  sum_disc_price_inst_cmd_firstIdx        <= l_sum_disc_price_cmd_firstIdx;
  sum_disc_price_inst_cmd_lastIdx         <= l_sum_disc_price_cmd_lastIdx;
  sum_disc_price_inst_cmd_ctrl            <= l_sum_disc_price_cmd_ctrl;
  sum_disc_price_inst_cmd_tag             <= l_sum_disc_price_cmd_tag;

  sum_disc_price_inst_in_valid(0)         <= l_sum_disc_price_valid;
  l_sum_disc_price_ready                  <= sum_disc_price_inst_in_ready(0);
  sum_disc_price_inst_in_data             <= l_sum_disc_price;
  sum_disc_price_inst_in_dvalid(0)        <= l_sum_disc_price_dvalid;
  sum_disc_price_inst_in_last(0)          <= l_sum_disc_price_last;

  sum_charge_inst_cmd_valid               <= l_sum_charge_cmd_valid;
  l_sum_charge_cmd_ready                  <= sum_charge_inst_cmd_ready;
  sum_charge_inst_cmd_firstIdx            <= l_sum_charge_cmd_firstIdx;
  sum_charge_inst_cmd_lastIdx             <= l_sum_charge_cmd_lastIdx;
  sum_charge_inst_cmd_ctrl                <= l_sum_charge_cmd_ctrl;
  sum_charge_inst_cmd_tag                 <= l_sum_charge_cmd_tag;

  sum_charge_inst_in_valid(0)             <= l_sum_charge_valid;
  l_sum_charge_ready                      <= sum_charge_inst_in_ready(0);
  sum_charge_inst_in_data                 <= l_sum_charge;
  sum_charge_inst_in_dvalid(0)            <= l_sum_charge_dvalid;
  sum_charge_inst_in_last(0)              <= l_sum_charge_last;

  avg_qty_inst_cmd_valid                  <= l_avg_qty_cmd_valid;
  l_avg_qty_cmd_ready                     <= avg_qty_inst_cmd_ready;
  avg_qty_inst_cmd_firstIdx               <= l_avg_qty_cmd_firstIdx;
  avg_qty_inst_cmd_lastIdx                <= l_avg_qty_cmd_lastIdx;
  avg_qty_inst_cmd_ctrl                   <= l_avg_qty_cmd_ctrl;
  avg_qty_inst_cmd_tag                    <= l_avg_qty_cmd_tag;

  avg_qty_inst_in_valid(0)                <= l_avg_qty_valid;
  l_avg_qty_ready                         <= avg_qty_inst_in_ready(0);
  avg_qty_inst_in_data                    <= l_avg_qty;
  avg_qty_inst_in_dvalid(0)               <= l_avg_qty_dvalid;
  avg_qty_inst_in_last(0)                 <= l_avg_qty_last;

  avg_price_inst_cmd_valid                <= l_avg_price_cmd_valid;
  l_avg_price_cmd_ready                   <= avg_price_inst_cmd_ready;
  avg_price_inst_cmd_firstIdx             <= l_avg_price_cmd_firstIdx;
  avg_price_inst_cmd_lastIdx              <= l_avg_price_cmd_lastIdx;
  avg_price_inst_cmd_ctrl                 <= l_avg_price_cmd_ctrl;
  avg_price_inst_cmd_tag                  <= l_avg_price_cmd_tag;

  avg_price_inst_in_valid(0)              <= l_avg_price_valid;
  l_avg_price_ready                       <= avg_price_inst_in_ready(0);
  avg_price_inst_in_data                  <= l_avg_price;
  avg_price_inst_in_dvalid(0)             <= l_avg_price_dvalid;
  avg_price_inst_in_last(0)               <= l_avg_price_last;

  avg_disc_inst_cmd_valid                 <= l_avg_disc_cmd_valid;
  l_avg_disc_cmd_ready                    <= avg_disc_inst_cmd_ready;
  avg_disc_inst_cmd_firstIdx              <= l_avg_disc_cmd_firstIdx;
  avg_disc_inst_cmd_lastIdx               <= l_avg_disc_cmd_lastIdx;
  avg_disc_inst_cmd_ctrl                  <= l_avg_disc_cmd_ctrl;
  avg_disc_inst_cmd_tag                   <= l_avg_disc_cmd_tag;

  avg_disc_inst_in_valid(0)               <= l_avg_disc_valid;
  l_avg_disc_ready                        <= avg_disc_inst_in_ready(0);
  avg_disc_inst_in_data                   <= l_avg_disc;
  avg_disc_inst_in_dvalid(0)              <= l_avg_disc_dvalid;
  avg_disc_inst_in_last(0)                <= l_avg_disc_last;

  count_order_inst_cmd_valid              <= l_count_order_cmd_valid;
  l_count_order_cmd_ready                 <= count_order_inst_cmd_ready;
  count_order_inst_cmd_firstIdx           <= l_count_order_cmd_firstIdx;
  count_order_inst_cmd_lastIdx            <= l_count_order_cmd_lastIdx;
  count_order_inst_cmd_ctrl               <= l_count_order_cmd_ctrl;
  count_order_inst_cmd_tag                <= l_count_order_cmd_tag;

  count_order_inst_in_valid(0)            <= l_count_order_valid;
  l_count_order_ready                     <= count_order_inst_in_ready(0);
  count_order_inst_in_data                <= l_count_order;
  count_order_inst_in_dvalid(0)           <= l_count_order_dvalid;
  count_order_inst_in_last(0)             <= l_count_order_last;

  quantity_inst : ArrayReader
  generic map(
    BUS_ADDR_WIDTH     => L_QUANTITY_BUS_ADDR_WIDTH,
    BUS_DATA_WIDTH     => L_QUANTITY_BUS_DATA_WIDTH,
    BUS_LEN_WIDTH      => L_QUANTITY_BUS_LEN_WIDTH,
    BUS_BURST_STEP_LEN => L_QUANTITY_BUS_BURST_STEP_LEN,
    BUS_BURST_MAX_LEN  => L_QUANTITY_BUS_BURST_MAX_LEN,
    INDEX_WIDTH        => INDEX_WIDTH,
    CFG                => "prim(64)",
    CMD_TAG_ENABLE     => true,
    CMD_TAG_WIDTH      => TAG_WIDTH
  )
  port map(
    bcd_clk        => bcd_clk,
    bcd_reset      => bcd_reset,
    kcd_clk        => kcd_clk,
    kcd_reset      => kcd_reset,
    cmd_valid      => quantity_inst_cmd_valid,
    cmd_ready      => quantity_inst_cmd_ready,
    cmd_firstIdx   => quantity_inst_cmd_firstIdx,
    cmd_lastIdx    => quantity_inst_cmd_lastIdx,
    cmd_ctrl       => quantity_inst_cmd_ctrl,
    cmd_tag        => quantity_inst_cmd_tag,
    unl_valid      => quantity_inst_unl_valid,
    unl_ready      => quantity_inst_unl_ready,
    unl_tag        => quantity_inst_unl_tag,
    bus_rreq_valid => quantity_inst_bus_rreq_valid,
    bus_rreq_ready => quantity_inst_bus_rreq_ready,
    bus_rreq_addr  => quantity_inst_bus_rreq_addr,
    bus_rreq_len   => quantity_inst_bus_rreq_len,
    bus_rdat_valid => quantity_inst_bus_rdat_valid,
    bus_rdat_ready => quantity_inst_bus_rdat_ready,
    bus_rdat_data  => quantity_inst_bus_rdat_data,
    bus_rdat_last  => quantity_inst_bus_rdat_last,
    out_valid      => quantity_inst_out_valid,
    out_ready      => quantity_inst_out_ready,
    out_data       => quantity_inst_out_data,
    out_dvalid     => quantity_inst_out_dvalid,
    out_last       => quantity_inst_out_last
  );

  extendedprice_inst : ArrayReader
  generic map(
    BUS_ADDR_WIDTH     => L_EXTENDEDPRICE_BUS_ADDR_WIDTH,
    BUS_DATA_WIDTH     => L_EXTENDEDPRICE_BUS_DATA_WIDTH,
    BUS_LEN_WIDTH      => L_EXTENDEDPRICE_BUS_LEN_WIDTH,
    BUS_BURST_STEP_LEN => L_EXTENDEDPRICE_BUS_BURST_STEP_LEN,
    BUS_BURST_MAX_LEN  => L_EXTENDEDPRICE_BUS_BURST_MAX_LEN,
    INDEX_WIDTH        => INDEX_WIDTH,
    CFG                => "prim(64)",
    CMD_TAG_ENABLE     => true,
    CMD_TAG_WIDTH      => TAG_WIDTH
  )
  port map(
    bcd_clk        => bcd_clk,
    bcd_reset      => bcd_reset,
    kcd_clk        => kcd_clk,
    kcd_reset      => kcd_reset,
    cmd_valid      => extendedprice_inst_cmd_valid,
    cmd_ready      => extendedprice_inst_cmd_ready,
    cmd_firstIdx   => extendedprice_inst_cmd_firstIdx,
    cmd_lastIdx    => extendedprice_inst_cmd_lastIdx,
    cmd_ctrl       => extendedprice_inst_cmd_ctrl,
    cmd_tag        => extendedprice_inst_cmd_tag,
    unl_valid      => extendedprice_inst_unl_valid,
    unl_ready      => extendedprice_inst_unl_ready,
    unl_tag        => extendedprice_inst_unl_tag,
    bus_rreq_valid => extendedprice_inst_bus_rreq_valid,
    bus_rreq_ready => extendedprice_inst_bus_rreq_ready,
    bus_rreq_addr  => extendedprice_inst_bus_rreq_addr,
    bus_rreq_len   => extendedprice_inst_bus_rreq_len,
    bus_rdat_valid => extendedprice_inst_bus_rdat_valid,
    bus_rdat_ready => extendedprice_inst_bus_rdat_ready,
    bus_rdat_data  => extendedprice_inst_bus_rdat_data,
    bus_rdat_last  => extendedprice_inst_bus_rdat_last,
    out_valid      => extendedprice_inst_out_valid,
    out_ready      => extendedprice_inst_out_ready,
    out_data       => extendedprice_inst_out_data,
    out_dvalid     => extendedprice_inst_out_dvalid,
    out_last       => extendedprice_inst_out_last
  );

  discount_inst : ArrayReader
  generic map(
    BUS_ADDR_WIDTH     => L_DISCOUNT_BUS_ADDR_WIDTH,
    BUS_DATA_WIDTH     => L_DISCOUNT_BUS_DATA_WIDTH,
    BUS_LEN_WIDTH      => L_DISCOUNT_BUS_LEN_WIDTH,
    BUS_BURST_STEP_LEN => L_DISCOUNT_BUS_BURST_STEP_LEN,
    BUS_BURST_MAX_LEN  => L_DISCOUNT_BUS_BURST_MAX_LEN,
    INDEX_WIDTH        => INDEX_WIDTH,
    CFG                => "prim(64)",
    CMD_TAG_ENABLE     => true,
    CMD_TAG_WIDTH      => TAG_WIDTH
  )
  port map(
    bcd_clk        => bcd_clk,
    bcd_reset      => bcd_reset,
    kcd_clk        => kcd_clk,
    kcd_reset      => kcd_reset,
    cmd_valid      => discount_inst_cmd_valid,
    cmd_ready      => discount_inst_cmd_ready,
    cmd_firstIdx   => discount_inst_cmd_firstIdx,
    cmd_lastIdx    => discount_inst_cmd_lastIdx,
    cmd_ctrl       => discount_inst_cmd_ctrl,
    cmd_tag        => discount_inst_cmd_tag,
    unl_valid      => discount_inst_unl_valid,
    unl_ready      => discount_inst_unl_ready,
    unl_tag        => discount_inst_unl_tag,
    bus_rreq_valid => discount_inst_bus_rreq_valid,
    bus_rreq_ready => discount_inst_bus_rreq_ready,
    bus_rreq_addr  => discount_inst_bus_rreq_addr,
    bus_rreq_len   => discount_inst_bus_rreq_len,
    bus_rdat_valid => discount_inst_bus_rdat_valid,
    bus_rdat_ready => discount_inst_bus_rdat_ready,
    bus_rdat_data  => discount_inst_bus_rdat_data,
    bus_rdat_last  => discount_inst_bus_rdat_last,
    out_valid      => discount_inst_out_valid,
    out_ready      => discount_inst_out_ready,
    out_data       => discount_inst_out_data,
    out_dvalid     => discount_inst_out_dvalid,
    out_last       => discount_inst_out_last
  );

  tax_inst : ArrayReader
  generic map(
    BUS_ADDR_WIDTH     => L_TAX_BUS_ADDR_WIDTH,
    BUS_DATA_WIDTH     => L_TAX_BUS_DATA_WIDTH,
    BUS_LEN_WIDTH      => L_TAX_BUS_LEN_WIDTH,
    BUS_BURST_STEP_LEN => L_TAX_BUS_BURST_STEP_LEN,
    BUS_BURST_MAX_LEN  => L_TAX_BUS_BURST_MAX_LEN,
    INDEX_WIDTH        => INDEX_WIDTH,
    CFG                => "prim(64)",
    CMD_TAG_ENABLE     => true,
    CMD_TAG_WIDTH      => TAG_WIDTH
  )
  port map(
    bcd_clk        => bcd_clk,
    bcd_reset      => bcd_reset,
    kcd_clk        => kcd_clk,
    kcd_reset      => kcd_reset,
    cmd_valid      => tax_inst_cmd_valid,
    cmd_ready      => tax_inst_cmd_ready,
    cmd_firstIdx   => tax_inst_cmd_firstIdx,
    cmd_lastIdx    => tax_inst_cmd_lastIdx,
    cmd_ctrl       => tax_inst_cmd_ctrl,
    cmd_tag        => tax_inst_cmd_tag,
    unl_valid      => tax_inst_unl_valid,
    unl_ready      => tax_inst_unl_ready,
    unl_tag        => tax_inst_unl_tag,
    bus_rreq_valid => tax_inst_bus_rreq_valid,
    bus_rreq_ready => tax_inst_bus_rreq_ready,
    bus_rreq_addr  => tax_inst_bus_rreq_addr,
    bus_rreq_len   => tax_inst_bus_rreq_len,
    bus_rdat_valid => tax_inst_bus_rdat_valid,
    bus_rdat_ready => tax_inst_bus_rdat_ready,
    bus_rdat_data  => tax_inst_bus_rdat_data,
    bus_rdat_last  => tax_inst_bus_rdat_last,
    out_valid      => tax_inst_out_valid,
    out_ready      => tax_inst_out_ready,
    out_data       => tax_inst_out_data,
    out_dvalid     => tax_inst_out_dvalid,
    out_last       => tax_inst_out_last
  );

  returnflag_inst : ArrayReader
  generic map(
    BUS_ADDR_WIDTH     => L_RETURNFLAG_BUS_ADDR_WIDTH,
    BUS_DATA_WIDTH     => L_RETURNFLAG_BUS_DATA_WIDTH,
    BUS_LEN_WIDTH      => L_RETURNFLAG_BUS_LEN_WIDTH,
    BUS_BURST_STEP_LEN => L_RETURNFLAG_BUS_BURST_STEP_LEN,
    BUS_BURST_MAX_LEN  => L_RETURNFLAG_BUS_BURST_MAX_LEN,
    INDEX_WIDTH        => INDEX_WIDTH,
    CFG                => "listprim(8)",
    CMD_TAG_ENABLE     => true,
    CMD_TAG_WIDTH      => TAG_WIDTH
  )
  port map(
    bcd_clk        => bcd_clk,
    bcd_reset      => bcd_reset,
    kcd_clk        => kcd_clk,
    kcd_reset      => kcd_reset,
    cmd_valid      => returnflag_inst_cmd_valid,
    cmd_ready      => returnflag_inst_cmd_ready,
    cmd_firstIdx   => returnflag_inst_cmd_firstIdx,
    cmd_lastIdx    => returnflag_inst_cmd_lastIdx,
    cmd_ctrl       => returnflag_inst_cmd_ctrl,
    cmd_tag        => returnflag_inst_cmd_tag,
    unl_valid      => returnflag_inst_unl_valid,
    unl_ready      => returnflag_inst_unl_ready,
    unl_tag        => returnflag_inst_unl_tag,
    bus_rreq_valid => returnflag_inst_bus_rreq_valid,
    bus_rreq_ready => returnflag_inst_bus_rreq_ready,
    bus_rreq_addr  => returnflag_inst_bus_rreq_addr,
    bus_rreq_len   => returnflag_inst_bus_rreq_len,
    bus_rdat_valid => returnflag_inst_bus_rdat_valid,
    bus_rdat_ready => returnflag_inst_bus_rdat_ready,
    bus_rdat_data  => returnflag_inst_bus_rdat_data,
    bus_rdat_last  => returnflag_inst_bus_rdat_last,
    out_valid      => returnflag_inst_out_valid,
    out_ready      => returnflag_inst_out_ready,
    out_data       => returnflag_inst_out_data,
    out_dvalid     => returnflag_inst_out_dvalid,
    out_last       => returnflag_inst_out_last
  );

  linestatus_inst : ArrayReader
  generic map(
    BUS_ADDR_WIDTH     => L_LINESTATUS_BUS_ADDR_WIDTH,
    BUS_DATA_WIDTH     => L_LINESTATUS_BUS_DATA_WIDTH,
    BUS_LEN_WIDTH      => L_LINESTATUS_BUS_LEN_WIDTH,
    BUS_BURST_STEP_LEN => L_LINESTATUS_BUS_BURST_STEP_LEN,
    BUS_BURST_MAX_LEN  => L_LINESTATUS_BUS_BURST_MAX_LEN,
    INDEX_WIDTH        => INDEX_WIDTH,
    CFG                => "listprim(8)",
    CMD_TAG_ENABLE     => true,
    CMD_TAG_WIDTH      => TAG_WIDTH
  )
  port map(
    bcd_clk        => bcd_clk,
    bcd_reset      => bcd_reset,
    kcd_clk        => kcd_clk,
    kcd_reset      => kcd_reset,
    cmd_valid      => linestatus_inst_cmd_valid,
    cmd_ready      => linestatus_inst_cmd_ready,
    cmd_firstIdx   => linestatus_inst_cmd_firstIdx,
    cmd_lastIdx    => linestatus_inst_cmd_lastIdx,
    cmd_ctrl       => linestatus_inst_cmd_ctrl,
    cmd_tag        => linestatus_inst_cmd_tag,
    unl_valid      => linestatus_inst_unl_valid,
    unl_ready      => linestatus_inst_unl_ready,
    unl_tag        => linestatus_inst_unl_tag,
    bus_rreq_valid => linestatus_inst_bus_rreq_valid,
    bus_rreq_ready => linestatus_inst_bus_rreq_ready,
    bus_rreq_addr  => linestatus_inst_bus_rreq_addr,
    bus_rreq_len   => linestatus_inst_bus_rreq_len,
    bus_rdat_valid => linestatus_inst_bus_rdat_valid,
    bus_rdat_ready => linestatus_inst_bus_rdat_ready,
    bus_rdat_data  => linestatus_inst_bus_rdat_data,
    bus_rdat_last  => linestatus_inst_bus_rdat_last,
    out_valid      => linestatus_inst_out_valid,
    out_ready      => linestatus_inst_out_ready,
    out_data       => linestatus_inst_out_data,
    out_dvalid     => linestatus_inst_out_dvalid,
    out_last       => linestatus_inst_out_last
  );

  shipdate_inst : ArrayReader
  generic map(
    BUS_ADDR_WIDTH     => L_SHIPDATE_BUS_ADDR_WIDTH,
    BUS_DATA_WIDTH     => L_SHIPDATE_BUS_DATA_WIDTH,
    BUS_LEN_WIDTH      => L_SHIPDATE_BUS_LEN_WIDTH,
    BUS_BURST_STEP_LEN => L_SHIPDATE_BUS_BURST_STEP_LEN,
    BUS_BURST_MAX_LEN  => L_SHIPDATE_BUS_BURST_MAX_LEN,
    INDEX_WIDTH        => INDEX_WIDTH,
    CFG                => "prim(32)",
    CMD_TAG_ENABLE     => true,
    CMD_TAG_WIDTH      => TAG_WIDTH
  )
  port map(
    bcd_clk        => bcd_clk,
    bcd_reset      => bcd_reset,
    kcd_clk        => kcd_clk,
    kcd_reset      => kcd_reset,
    cmd_valid      => shipdate_inst_cmd_valid,
    cmd_ready      => shipdate_inst_cmd_ready,
    cmd_firstIdx   => shipdate_inst_cmd_firstIdx,
    cmd_lastIdx    => shipdate_inst_cmd_lastIdx,
    cmd_ctrl       => shipdate_inst_cmd_ctrl,
    cmd_tag        => shipdate_inst_cmd_tag,
    unl_valid      => shipdate_inst_unl_valid,
    unl_ready      => shipdate_inst_unl_ready,
    unl_tag        => shipdate_inst_unl_tag,
    bus_rreq_valid => shipdate_inst_bus_rreq_valid,
    bus_rreq_ready => shipdate_inst_bus_rreq_ready,
    bus_rreq_addr  => shipdate_inst_bus_rreq_addr,
    bus_rreq_len   => shipdate_inst_bus_rreq_len,
    bus_rdat_valid => shipdate_inst_bus_rdat_valid,
    bus_rdat_ready => shipdate_inst_bus_rdat_ready,
    bus_rdat_data  => shipdate_inst_bus_rdat_data,
    bus_rdat_last  => shipdate_inst_bus_rdat_last,
    out_valid      => shipdate_inst_out_valid,
    out_ready      => shipdate_inst_out_ready,
    out_data       => shipdate_inst_out_data,
    out_dvalid     => shipdate_inst_out_dvalid,
    out_last       => shipdate_inst_out_last
  );

  l_quantity_valid                  <= quantity_inst_out_valid(0);
  quantity_inst_out_ready(0)        <= l_quantity_ready;
  l_quantity_dvalid                 <= quantity_inst_out_dvalid(0);
  l_quantity_last                   <= quantity_inst_out_last(0);
  l_quantity                        <= quantity_inst_out_data;

  l_quantity_bus_rreq_valid         <= quantity_inst_bus_rreq_valid;
  quantity_inst_bus_rreq_ready      <= l_quantity_bus_rreq_ready;
  l_quantity_bus_rreq_addr          <= quantity_inst_bus_rreq_addr;
  l_quantity_bus_rreq_len           <= quantity_inst_bus_rreq_len;
  quantity_inst_bus_rdat_valid      <= l_quantity_bus_rdat_valid;
  l_quantity_bus_rdat_ready         <= quantity_inst_bus_rdat_ready;
  quantity_inst_bus_rdat_data       <= l_quantity_bus_rdat_data;
  quantity_inst_bus_rdat_last       <= l_quantity_bus_rdat_last;

  l_quantity_unl_valid              <= quantity_inst_unl_valid;
  quantity_inst_unl_ready           <= l_quantity_unl_ready;
  l_quantity_unl_tag                <= quantity_inst_unl_tag;

  l_extendedprice_valid             <= extendedprice_inst_out_valid(0);
  extendedprice_inst_out_ready(0)   <= l_extendedprice_ready;
  l_extendedprice_dvalid            <= extendedprice_inst_out_dvalid(0);
  l_extendedprice_last              <= extendedprice_inst_out_last(0);
  l_extendedprice                   <= extendedprice_inst_out_data;

  l_extendedprice_bus_rreq_valid    <= extendedprice_inst_bus_rreq_valid;
  extendedprice_inst_bus_rreq_ready <= l_extendedprice_bus_rreq_ready;
  l_extendedprice_bus_rreq_addr     <= extendedprice_inst_bus_rreq_addr;
  l_extendedprice_bus_rreq_len      <= extendedprice_inst_bus_rreq_len;
  extendedprice_inst_bus_rdat_valid <= l_extendedprice_bus_rdat_valid;
  l_extendedprice_bus_rdat_ready    <= extendedprice_inst_bus_rdat_ready;
  extendedprice_inst_bus_rdat_data  <= l_extendedprice_bus_rdat_data;
  extendedprice_inst_bus_rdat_last  <= l_extendedprice_bus_rdat_last;

  l_extendedprice_unl_valid         <= extendedprice_inst_unl_valid;
  extendedprice_inst_unl_ready      <= l_extendedprice_unl_ready;
  l_extendedprice_unl_tag           <= extendedprice_inst_unl_tag;

  l_discount_valid                  <= discount_inst_out_valid(0);
  discount_inst_out_ready(0)        <= l_discount_ready;
  l_discount_dvalid                 <= discount_inst_out_dvalid(0);
  l_discount_last                   <= discount_inst_out_last(0);
  l_discount                        <= discount_inst_out_data;

  l_discount_bus_rreq_valid         <= discount_inst_bus_rreq_valid;
  discount_inst_bus_rreq_ready      <= l_discount_bus_rreq_ready;
  l_discount_bus_rreq_addr          <= discount_inst_bus_rreq_addr;
  l_discount_bus_rreq_len           <= discount_inst_bus_rreq_len;
  discount_inst_bus_rdat_valid      <= l_discount_bus_rdat_valid;
  l_discount_bus_rdat_ready         <= discount_inst_bus_rdat_ready;
  discount_inst_bus_rdat_data       <= l_discount_bus_rdat_data;
  discount_inst_bus_rdat_last       <= l_discount_bus_rdat_last;

  l_discount_unl_valid              <= discount_inst_unl_valid;
  discount_inst_unl_ready           <= l_discount_unl_ready;
  l_discount_unl_tag                <= discount_inst_unl_tag;

  l_tax_valid                       <= tax_inst_out_valid(0);
  tax_inst_out_ready(0)             <= l_tax_ready;
  l_tax_dvalid                      <= tax_inst_out_dvalid(0);
  l_tax_last                        <= tax_inst_out_last(0);
  l_tax                             <= tax_inst_out_data;

  l_tax_bus_rreq_valid              <= tax_inst_bus_rreq_valid;
  tax_inst_bus_rreq_ready           <= l_tax_bus_rreq_ready;
  l_tax_bus_rreq_addr               <= tax_inst_bus_rreq_addr;
  l_tax_bus_rreq_len                <= tax_inst_bus_rreq_len;
  tax_inst_bus_rdat_valid           <= l_tax_bus_rdat_valid;
  l_tax_bus_rdat_ready              <= tax_inst_bus_rdat_ready;
  tax_inst_bus_rdat_data            <= l_tax_bus_rdat_data;
  tax_inst_bus_rdat_last            <= l_tax_bus_rdat_last;

  l_tax_unl_valid                   <= tax_inst_unl_valid;
  tax_inst_unl_ready                <= l_tax_unl_ready;
  l_tax_unl_tag                     <= tax_inst_unl_tag;

  l_returnflag_valid                <= returnflag_inst_out_valid(0);
  l_returnflag_chars_valid          <= returnflag_inst_out_valid(1);
  returnflag_inst_out_ready(0)      <= l_returnflag_ready;
  returnflag_inst_out_ready(1)      <= l_returnflag_chars_ready;
  l_returnflag_dvalid               <= returnflag_inst_out_dvalid(0);
  l_returnflag_chars_dvalid         <= returnflag_inst_out_dvalid(1);
  l_returnflag_last                 <= returnflag_inst_out_last(0);
  l_returnflag_chars_last           <= returnflag_inst_out_last(1);
  l_returnflag_length               <= returnflag_inst_out_data(31 downto 0);
  l_returnflag_count                <= returnflag_inst_out_data(32 downto 32);
  l_returnflag_chars                <= returnflag_inst_out_data(40 downto 33);
  l_returnflag_chars_count          <= returnflag_inst_out_data(41 downto 41);

  l_returnflag_bus_rreq_valid       <= returnflag_inst_bus_rreq_valid;
  returnflag_inst_bus_rreq_ready    <= l_returnflag_bus_rreq_ready;
  l_returnflag_bus_rreq_addr        <= returnflag_inst_bus_rreq_addr;
  l_returnflag_bus_rreq_len         <= returnflag_inst_bus_rreq_len;
  returnflag_inst_bus_rdat_valid    <= l_returnflag_bus_rdat_valid;
  l_returnflag_bus_rdat_ready       <= returnflag_inst_bus_rdat_ready;
  returnflag_inst_bus_rdat_data     <= l_returnflag_bus_rdat_data;
  returnflag_inst_bus_rdat_last     <= l_returnflag_bus_rdat_last;

  l_returnflag_unl_valid            <= returnflag_inst_unl_valid;
  returnflag_inst_unl_ready         <= l_returnflag_unl_ready;
  l_returnflag_unl_tag              <= returnflag_inst_unl_tag;

  l_linestatus_valid                <= linestatus_inst_out_valid(0);
  l_linestatus_chars_valid          <= linestatus_inst_out_valid(1);
  linestatus_inst_out_ready(0)      <= l_linestatus_ready;
  linestatus_inst_out_ready(1)      <= l_linestatus_chars_ready;
  l_linestatus_dvalid               <= linestatus_inst_out_dvalid(0);
  l_linestatus_chars_dvalid         <= linestatus_inst_out_dvalid(1);
  l_linestatus_last                 <= linestatus_inst_out_last(0);
  l_linestatus_chars_last           <= linestatus_inst_out_last(1);
  l_linestatus_length               <= linestatus_inst_out_data(31 downto 0);
  l_linestatus_count                <= linestatus_inst_out_data(32 downto 32);
  l_linestatus_chars                <= linestatus_inst_out_data(40 downto 33);
  l_linestatus_chars_count          <= linestatus_inst_out_data(41 downto 41);

  l_linestatus_bus_rreq_valid       <= linestatus_inst_bus_rreq_valid;
  linestatus_inst_bus_rreq_ready    <= l_linestatus_bus_rreq_ready;
  l_linestatus_bus_rreq_addr        <= linestatus_inst_bus_rreq_addr;
  l_linestatus_bus_rreq_len         <= linestatus_inst_bus_rreq_len;
  linestatus_inst_bus_rdat_valid    <= l_linestatus_bus_rdat_valid;
  l_linestatus_bus_rdat_ready       <= linestatus_inst_bus_rdat_ready;
  linestatus_inst_bus_rdat_data     <= l_linestatus_bus_rdat_data;
  linestatus_inst_bus_rdat_last     <= l_linestatus_bus_rdat_last;

  l_linestatus_unl_valid            <= linestatus_inst_unl_valid;
  linestatus_inst_unl_ready         <= l_linestatus_unl_ready;
  l_linestatus_unl_tag              <= linestatus_inst_unl_tag;

  l_shipdate_valid                  <= shipdate_inst_out_valid(0);
  shipdate_inst_out_ready(0)        <= l_shipdate_ready;
  l_shipdate_dvalid                 <= shipdate_inst_out_dvalid(0);
  l_shipdate_last                   <= shipdate_inst_out_last(0);
  l_shipdate                        <= shipdate_inst_out_data;

  l_shipdate_bus_rreq_valid         <= shipdate_inst_bus_rreq_valid;
  shipdate_inst_bus_rreq_ready      <= l_shipdate_bus_rreq_ready;
  l_shipdate_bus_rreq_addr          <= shipdate_inst_bus_rreq_addr;
  l_shipdate_bus_rreq_len           <= shipdate_inst_bus_rreq_len;
  shipdate_inst_bus_rdat_valid      <= l_shipdate_bus_rdat_valid;
  l_shipdate_bus_rdat_ready         <= shipdate_inst_bus_rdat_ready;
  shipdate_inst_bus_rdat_data       <= l_shipdate_bus_rdat_data;
  shipdate_inst_bus_rdat_last       <= l_shipdate_bus_rdat_last;

  l_shipdate_unl_valid              <= shipdate_inst_unl_valid;
  shipdate_inst_unl_ready           <= l_shipdate_unl_ready;
  l_shipdate_unl_tag                <= shipdate_inst_unl_tag;

  quantity_inst_cmd_valid           <= l_quantity_cmd_valid;
  l_quantity_cmd_ready              <= quantity_inst_cmd_ready;
  quantity_inst_cmd_firstIdx        <= l_quantity_cmd_firstIdx;
  quantity_inst_cmd_lastIdx         <= l_quantity_cmd_lastIdx;
  quantity_inst_cmd_ctrl            <= l_quantity_cmd_ctrl;
  quantity_inst_cmd_tag             <= l_quantity_cmd_tag;

  extendedprice_inst_cmd_valid      <= l_extendedprice_cmd_valid;
  l_extendedprice_cmd_ready         <= extendedprice_inst_cmd_ready;
  extendedprice_inst_cmd_firstIdx   <= l_extendedprice_cmd_firstIdx;
  extendedprice_inst_cmd_lastIdx    <= l_extendedprice_cmd_lastIdx;
  extendedprice_inst_cmd_ctrl       <= l_extendedprice_cmd_ctrl;
  extendedprice_inst_cmd_tag        <= l_extendedprice_cmd_tag;

  discount_inst_cmd_valid           <= l_discount_cmd_valid;
  l_discount_cmd_ready              <= discount_inst_cmd_ready;
  discount_inst_cmd_firstIdx        <= l_discount_cmd_firstIdx;
  discount_inst_cmd_lastIdx         <= l_discount_cmd_lastIdx;
  discount_inst_cmd_ctrl            <= l_discount_cmd_ctrl;
  discount_inst_cmd_tag             <= l_discount_cmd_tag;

  tax_inst_cmd_valid                <= l_tax_cmd_valid;
  l_tax_cmd_ready                   <= tax_inst_cmd_ready;
  tax_inst_cmd_firstIdx             <= l_tax_cmd_firstIdx;
  tax_inst_cmd_lastIdx              <= l_tax_cmd_lastIdx;
  tax_inst_cmd_ctrl                 <= l_tax_cmd_ctrl;
  tax_inst_cmd_tag                  <= l_tax_cmd_tag;

  returnflag_inst_cmd_valid         <= l_returnflag_cmd_valid;
  l_returnflag_cmd_ready            <= returnflag_inst_cmd_ready;
  returnflag_inst_cmd_firstIdx      <= l_returnflag_cmd_firstIdx;
  returnflag_inst_cmd_lastIdx       <= l_returnflag_cmd_lastIdx;
  returnflag_inst_cmd_ctrl          <= l_returnflag_cmd_ctrl;
  returnflag_inst_cmd_tag           <= l_returnflag_cmd_tag;

  linestatus_inst_cmd_valid         <= l_linestatus_cmd_valid;
  l_linestatus_cmd_ready            <= linestatus_inst_cmd_ready;
  linestatus_inst_cmd_firstIdx      <= l_linestatus_cmd_firstIdx;
  linestatus_inst_cmd_lastIdx       <= l_linestatus_cmd_lastIdx;
  linestatus_inst_cmd_ctrl          <= l_linestatus_cmd_ctrl;
  linestatus_inst_cmd_tag           <= l_linestatus_cmd_tag;

  shipdate_inst_cmd_valid           <= l_shipdate_cmd_valid;
  l_shipdate_cmd_ready              <= shipdate_inst_cmd_ready;
  shipdate_inst_cmd_firstIdx        <= l_shipdate_cmd_firstIdx;
  shipdate_inst_cmd_lastIdx         <= l_shipdate_cmd_lastIdx;
  shipdate_inst_cmd_ctrl            <= l_shipdate_cmd_ctrl;
  shipdate_inst_cmd_tag             <= l_shipdate_cmd_tag;

end architecture;