-- Copyright 2018-2019 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
-- This file was generated by Fletchgen. Modify this file at your own risk.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.Interconnect_pkg.all;

entity PriceSummary_Mantle is
  generic (
    INDEX_WIDTH        : integer := 32;
    TAG_WIDTH          : integer := 1;
    BUS_ADDR_WIDTH     : integer := 64;
    BUS_DATA_WIDTH     : integer := 512;
    BUS_LEN_WIDTH      : integer := 8;
    BUS_BURST_STEP_LEN : integer := 1;
    BUS_BURST_MAX_LEN  : integer := 16
  );
  port (
    bcd_clk            : in std_logic;
    bcd_reset          : in std_logic;
    kcd_clk            : in std_logic;
    kcd_reset          : in std_logic;
    mmio_awvalid       : in std_logic;
    mmio_awready       : out std_logic;
    mmio_awaddr        : in std_logic_vector(31 downto 0);
    mmio_wvalid        : in std_logic;
    mmio_wready        : out std_logic;
    mmio_wdata         : in std_logic_vector(31 downto 0);
    mmio_wstrb         : in std_logic_vector(3 downto 0);
    mmio_bvalid        : out std_logic;
    mmio_bready        : in std_logic;
    mmio_bresp         : out std_logic_vector(1 downto 0);
    mmio_arvalid       : in std_logic;
    mmio_arready       : out std_logic;
    mmio_araddr        : in std_logic_vector(31 downto 0);
    mmio_rvalid        : out std_logic;
    mmio_rready        : in std_logic;
    mmio_rdata         : out std_logic_vector(31 downto 0);
    mmio_rresp         : out std_logic_vector(1 downto 0);
    rd_mst_rreq_valid  : out std_logic;
    rd_mst_rreq_ready  : in std_logic;
    rd_mst_rreq_addr   : out std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
    rd_mst_rreq_len    : out std_logic_vector(BUS_LEN_WIDTH - 1 downto 0);
    rd_mst_rdat_valid  : in std_logic;
    rd_mst_rdat_ready  : out std_logic;
    rd_mst_rdat_data   : in std_logic_vector(BUS_DATA_WIDTH - 1 downto 0);
    rd_mst_rdat_last   : in std_logic;
    wr_mst_wreq_valid  : out std_logic;
    wr_mst_wreq_ready  : in std_logic;
    wr_mst_wreq_addr   : out std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
    wr_mst_wreq_len    : out std_logic_vector(BUS_LEN_WIDTH - 1 downto 0);
    wr_mst_wdat_valid  : out std_logic;
    wr_mst_wdat_ready  : in std_logic;
    wr_mst_wdat_data   : out std_logic_vector(BUS_DATA_WIDTH - 1 downto 0);
    wr_mst_wdat_strobe : out std_logic_vector(BUS_DATA_WIDTH/8 - 1 downto 0);
    wr_mst_wdat_last   : out std_logic
  );
end entity;

architecture Implementation of PriceSummary_Mantle is
  component PriceSummary_Nucleus is
    generic (
      INDEX_WIDTH                     : integer := 32;
      TAG_WIDTH                       : integer := 1;
      L_QUANTITY_BUS_ADDR_WIDTH       : integer := 64;
      L_EXTENDEDPRICE_BUS_ADDR_WIDTH  : integer := 64;
      L_DISCOUNT_BUS_ADDR_WIDTH       : integer := 64;
      L_TAX_BUS_ADDR_WIDTH            : integer := 64;
      L_RETURNFLAG_BUS_ADDR_WIDTH     : integer := 64;
      L_LINESTATUS_BUS_ADDR_WIDTH     : integer := 64;
      L_SHIPDATE_BUS_ADDR_WIDTH       : integer := 64;
      L_RETURNFLAG_O_BUS_ADDR_WIDTH   : integer := 64;
      L_LINESTATUS_O_BUS_ADDR_WIDTH   : integer := 64;
      L_SUM_QTY_BUS_ADDR_WIDTH        : integer := 64;
      L_SUM_BASE_PRICE_BUS_ADDR_WIDTH : integer := 64;
      L_SUM_DISC_PRICE_BUS_ADDR_WIDTH : integer := 64;
      L_SUM_CHARGE_BUS_ADDR_WIDTH     : integer := 64;
      L_AVG_QTY_BUS_ADDR_WIDTH        : integer := 64;
      L_AVG_PRICE_BUS_ADDR_WIDTH      : integer := 64;
      L_AVG_DISC_BUS_ADDR_WIDTH       : integer := 64;
      L_COUNT_ORDER_BUS_ADDR_WIDTH    : integer := 64
    );
    port (
      kcd_clk                       : in std_logic;
      kcd_reset                     : in std_logic;
      mmio_awvalid                  : in std_logic;
      mmio_awready                  : out std_logic;
      mmio_awaddr                   : in std_logic_vector(31 downto 0);
      mmio_wvalid                   : in std_logic;
      mmio_wready                   : out std_logic;
      mmio_wdata                    : in std_logic_vector(31 downto 0);
      mmio_wstrb                    : in std_logic_vector(3 downto 0);
      mmio_bvalid                   : out std_logic;
      mmio_bready                   : in std_logic;
      mmio_bresp                    : out std_logic_vector(1 downto 0);
      mmio_arvalid                  : in std_logic;
      mmio_arready                  : out std_logic;
      mmio_araddr                   : in std_logic_vector(31 downto 0);
      mmio_rvalid                   : out std_logic;
      mmio_rready                   : in std_logic;
      mmio_rdata                    : out std_logic_vector(31 downto 0);
      mmio_rresp                    : out std_logic_vector(1 downto 0);
      l_quantity_valid              : in std_logic;
      l_quantity_ready              : out std_logic;
      l_quantity_dvalid             : in std_logic;
      l_quantity_last               : in std_logic;
      l_quantity                    : in std_logic_vector(63 downto 0);
      l_extendedprice_valid         : in std_logic;
      l_extendedprice_ready         : out std_logic;
      l_extendedprice_dvalid        : in std_logic;
      l_extendedprice_last          : in std_logic;
      l_extendedprice               : in std_logic_vector(63 downto 0);
      l_discount_valid              : in std_logic;
      l_discount_ready              : out std_logic;
      l_discount_dvalid             : in std_logic;
      l_discount_last               : in std_logic;
      l_discount                    : in std_logic_vector(63 downto 0);
      l_tax_valid                   : in std_logic;
      l_tax_ready                   : out std_logic;
      l_tax_dvalid                  : in std_logic;
      l_tax_last                    : in std_logic;
      l_tax                         : in std_logic_vector(63 downto 0);
      l_returnflag_valid            : in std_logic;
      l_returnflag_ready            : out std_logic;
      l_returnflag_dvalid           : in std_logic;
      l_returnflag_last             : in std_logic;
      l_returnflag_length           : in std_logic_vector(31 downto 0);
      l_returnflag_count            : in std_logic_vector(0 downto 0);
      l_returnflag_chars_valid      : in std_logic;
      l_returnflag_chars_ready      : out std_logic;
      l_returnflag_chars_dvalid     : in std_logic;
      l_returnflag_chars_last       : in std_logic;
      l_returnflag_chars            : in std_logic_vector(7 downto 0);
      l_returnflag_chars_count      : in std_logic_vector(0 downto 0);
      l_linestatus_valid            : in std_logic;
      l_linestatus_ready            : out std_logic;
      l_linestatus_dvalid           : in std_logic;
      l_linestatus_last             : in std_logic;
      l_linestatus_length           : in std_logic_vector(31 downto 0);
      l_linestatus_count            : in std_logic_vector(0 downto 0);
      l_linestatus_chars_valid      : in std_logic;
      l_linestatus_chars_ready      : out std_logic;
      l_linestatus_chars_dvalid     : in std_logic;
      l_linestatus_chars_last       : in std_logic;
      l_linestatus_chars            : in std_logic_vector(7 downto 0);
      l_linestatus_chars_count      : in std_logic_vector(0 downto 0);
      l_shipdate_valid              : in std_logic;
      l_shipdate_ready              : out std_logic;
      l_shipdate_dvalid             : in std_logic;
      l_shipdate_last               : in std_logic;
      l_shipdate                    : in std_logic_vector(31 downto 0);
      l_quantity_unl_valid          : in std_logic;
      l_quantity_unl_ready          : out std_logic;
      l_quantity_unl_tag            : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_extendedprice_unl_valid     : in std_logic;
      l_extendedprice_unl_ready     : out std_logic;
      l_extendedprice_unl_tag       : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_discount_unl_valid          : in std_logic;
      l_discount_unl_ready          : out std_logic;
      l_discount_unl_tag            : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_tax_unl_valid               : in std_logic;
      l_tax_unl_ready               : out std_logic;
      l_tax_unl_tag                 : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_returnflag_unl_valid        : in std_logic;
      l_returnflag_unl_ready        : out std_logic;
      l_returnflag_unl_tag          : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_linestatus_unl_valid        : in std_logic;
      l_linestatus_unl_ready        : out std_logic;
      l_linestatus_unl_tag          : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_shipdate_unl_valid          : in std_logic;
      l_shipdate_unl_ready          : out std_logic;
      l_shipdate_unl_tag            : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_quantity_cmd_valid          : out std_logic;
      l_quantity_cmd_ready          : in std_logic;
      l_quantity_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_quantity_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_quantity_cmd_ctrl           : out std_logic_vector(L_QUANTITY_BUS_ADDR_WIDTH - 1 downto 0);
      l_quantity_cmd_tag            : out std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_extendedprice_cmd_valid     : out std_logic;
      l_extendedprice_cmd_ready     : in std_logic;
      l_extendedprice_cmd_firstIdx  : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_extendedprice_cmd_lastIdx   : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_extendedprice_cmd_ctrl      : out std_logic_vector(L_EXTENDEDPRICE_BUS_ADDR_WIDTH - 1 downto 0);
      l_extendedprice_cmd_tag       : out std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_discount_cmd_valid          : out std_logic;
      l_discount_cmd_ready          : in std_logic;
      l_discount_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_discount_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_discount_cmd_ctrl           : out std_logic_vector(L_DISCOUNT_BUS_ADDR_WIDTH - 1 downto 0);
      l_discount_cmd_tag            : out std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_tax_cmd_valid               : out std_logic;
      l_tax_cmd_ready               : in std_logic;
      l_tax_cmd_firstIdx            : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_tax_cmd_lastIdx             : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_tax_cmd_ctrl                : out std_logic_vector(L_TAX_BUS_ADDR_WIDTH - 1 downto 0);
      l_tax_cmd_tag                 : out std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_returnflag_cmd_valid        : out std_logic;
      l_returnflag_cmd_ready        : in std_logic;
      l_returnflag_cmd_firstIdx     : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_returnflag_cmd_lastIdx      : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_returnflag_cmd_ctrl         : out std_logic_vector(L_RETURNFLAG_BUS_ADDR_WIDTH * 2 - 1 downto 0);
      l_returnflag_cmd_tag          : out std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_linestatus_cmd_valid        : out std_logic;
      l_linestatus_cmd_ready        : in std_logic;
      l_linestatus_cmd_firstIdx     : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_linestatus_cmd_lastIdx      : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_linestatus_cmd_ctrl         : out std_logic_vector(L_LINESTATUS_BUS_ADDR_WIDTH * 2 - 1 downto 0);
      l_linestatus_cmd_tag          : out std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_shipdate_cmd_valid          : out std_logic;
      l_shipdate_cmd_ready          : in std_logic;
      l_shipdate_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_shipdate_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_shipdate_cmd_ctrl           : out std_logic_vector(L_SHIPDATE_BUS_ADDR_WIDTH - 1 downto 0);
      l_shipdate_cmd_tag            : out std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_returnflag_o_valid          : out std_logic;
      l_returnflag_o_ready          : in std_logic;
      l_returnflag_o_dvalid         : out std_logic;
      l_returnflag_o_last           : out std_logic;
      l_returnflag_o_length         : out std_logic_vector(31 downto 0);
      l_returnflag_o_count          : out std_logic_vector(0 downto 0);
      l_returnflag_o_chars_valid    : out std_logic;
      l_returnflag_o_chars_ready    : in std_logic;
      l_returnflag_o_chars_dvalid   : out std_logic;
      l_returnflag_o_chars_last     : out std_logic;
      l_returnflag_o_chars          : out std_logic_vector(7 downto 0);
      l_returnflag_o_chars_count    : out std_logic_vector(0 downto 0);
      l_linestatus_o_valid          : out std_logic;
      l_linestatus_o_ready          : in std_logic;
      l_linestatus_o_dvalid         : out std_logic;
      l_linestatus_o_last           : out std_logic;
      l_linestatus_o_length         : out std_logic_vector(31 downto 0);
      l_linestatus_o_count          : out std_logic_vector(0 downto 0);
      l_linestatus_o_chars_valid    : out std_logic;
      l_linestatus_o_chars_ready    : in std_logic;
      l_linestatus_o_chars_dvalid   : out std_logic;
      l_linestatus_o_chars_last     : out std_logic;
      l_linestatus_o_chars          : out std_logic_vector(7 downto 0);
      l_linestatus_o_chars_count    : out std_logic_vector(0 downto 0);
      l_sum_qty_valid               : out std_logic;
      l_sum_qty_ready               : in std_logic;
      l_sum_qty_dvalid              : out std_logic;
      l_sum_qty_last                : out std_logic;
      l_sum_qty                     : out std_logic_vector(63 downto 0);
      l_sum_base_price_valid        : out std_logic;
      l_sum_base_price_ready        : in std_logic;
      l_sum_base_price_dvalid       : out std_logic;
      l_sum_base_price_last         : out std_logic;
      l_sum_base_price              : out std_logic_vector(63 downto 0);
      l_sum_disc_price_valid        : out std_logic;
      l_sum_disc_price_ready        : in std_logic;
      l_sum_disc_price_dvalid       : out std_logic;
      l_sum_disc_price_last         : out std_logic;
      l_sum_disc_price              : out std_logic_vector(63 downto 0);
      l_sum_charge_valid            : out std_logic;
      l_sum_charge_ready            : in std_logic;
      l_sum_charge_dvalid           : out std_logic;
      l_sum_charge_last             : out std_logic;
      l_sum_charge                  : out std_logic_vector(63 downto 0);
      l_avg_qty_valid               : out std_logic;
      l_avg_qty_ready               : in std_logic;
      l_avg_qty_dvalid              : out std_logic;
      l_avg_qty_last                : out std_logic;
      l_avg_qty                     : out std_logic_vector(63 downto 0);
      l_avg_price_valid             : out std_logic;
      l_avg_price_ready             : in std_logic;
      l_avg_price_dvalid            : out std_logic;
      l_avg_price_last              : out std_logic;
      l_avg_price                   : out std_logic_vector(63 downto 0);
      l_avg_disc_valid              : out std_logic;
      l_avg_disc_ready              : in std_logic;
      l_avg_disc_dvalid             : out std_logic;
      l_avg_disc_last               : out std_logic;
      l_avg_disc                    : out std_logic_vector(63 downto 0);
      l_count_order_valid           : out std_logic;
      l_count_order_ready           : in std_logic;
      l_count_order_dvalid          : out std_logic;
      l_count_order_last            : out std_logic;
      l_count_order                 : out std_logic_vector(63 downto 0);
      l_returnflag_o_unl_valid      : in std_logic;
      l_returnflag_o_unl_ready      : out std_logic;
      l_returnflag_o_unl_tag        : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_linestatus_o_unl_valid      : in std_logic;
      l_linestatus_o_unl_ready      : out std_logic;
      l_linestatus_o_unl_tag        : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_sum_qty_unl_valid           : in std_logic;
      l_sum_qty_unl_ready           : out std_logic;
      l_sum_qty_unl_tag             : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_sum_base_price_unl_valid    : in std_logic;
      l_sum_base_price_unl_ready    : out std_logic;
      l_sum_base_price_unl_tag      : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_sum_disc_price_unl_valid    : in std_logic;
      l_sum_disc_price_unl_ready    : out std_logic;
      l_sum_disc_price_unl_tag      : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_sum_charge_unl_valid        : in std_logic;
      l_sum_charge_unl_ready        : out std_logic;
      l_sum_charge_unl_tag          : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_avg_qty_unl_valid           : in std_logic;
      l_avg_qty_unl_ready           : out std_logic;
      l_avg_qty_unl_tag             : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_avg_price_unl_valid         : in std_logic;
      l_avg_price_unl_ready         : out std_logic;
      l_avg_price_unl_tag           : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_avg_disc_unl_valid          : in std_logic;
      l_avg_disc_unl_ready          : out std_logic;
      l_avg_disc_unl_tag            : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_count_order_unl_valid       : in std_logic;
      l_count_order_unl_ready       : out std_logic;
      l_count_order_unl_tag         : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_returnflag_o_cmd_valid      : out std_logic;
      l_returnflag_o_cmd_ready      : in std_logic;
      l_returnflag_o_cmd_firstIdx   : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_returnflag_o_cmd_lastIdx    : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_returnflag_o_cmd_ctrl       : out std_logic_vector(L_RETURNFLAG_O_BUS_ADDR_WIDTH * 2 - 1 downto 0);
      l_returnflag_o_cmd_tag        : out std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_linestatus_o_cmd_valid      : out std_logic;
      l_linestatus_o_cmd_ready      : in std_logic;
      l_linestatus_o_cmd_firstIdx   : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_linestatus_o_cmd_lastIdx    : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_linestatus_o_cmd_ctrl       : out std_logic_vector(L_LINESTATUS_O_BUS_ADDR_WIDTH * 2 - 1 downto 0);
      l_linestatus_o_cmd_tag        : out std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_sum_qty_cmd_valid           : out std_logic;
      l_sum_qty_cmd_ready           : in std_logic;
      l_sum_qty_cmd_firstIdx        : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_sum_qty_cmd_lastIdx         : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_sum_qty_cmd_ctrl            : out std_logic_vector(L_SUM_QTY_BUS_ADDR_WIDTH - 1 downto 0);
      l_sum_qty_cmd_tag             : out std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_sum_base_price_cmd_valid    : out std_logic;
      l_sum_base_price_cmd_ready    : in std_logic;
      l_sum_base_price_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_sum_base_price_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_sum_base_price_cmd_ctrl     : out std_logic_vector(L_SUM_BASE_PRICE_BUS_ADDR_WIDTH - 1 downto 0);
      l_sum_base_price_cmd_tag      : out std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_sum_disc_price_cmd_valid    : out std_logic;
      l_sum_disc_price_cmd_ready    : in std_logic;
      l_sum_disc_price_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_sum_disc_price_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_sum_disc_price_cmd_ctrl     : out std_logic_vector(L_SUM_DISC_PRICE_BUS_ADDR_WIDTH - 1 downto 0);
      l_sum_disc_price_cmd_tag      : out std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_sum_charge_cmd_valid        : out std_logic;
      l_sum_charge_cmd_ready        : in std_logic;
      l_sum_charge_cmd_firstIdx     : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_sum_charge_cmd_lastIdx      : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_sum_charge_cmd_ctrl         : out std_logic_vector(L_SUM_CHARGE_BUS_ADDR_WIDTH - 1 downto 0);
      l_sum_charge_cmd_tag          : out std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_avg_qty_cmd_valid           : out std_logic;
      l_avg_qty_cmd_ready           : in std_logic;
      l_avg_qty_cmd_firstIdx        : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_avg_qty_cmd_lastIdx         : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_avg_qty_cmd_ctrl            : out std_logic_vector(L_AVG_QTY_BUS_ADDR_WIDTH - 1 downto 0);
      l_avg_qty_cmd_tag             : out std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_avg_price_cmd_valid         : out std_logic;
      l_avg_price_cmd_ready         : in std_logic;
      l_avg_price_cmd_firstIdx      : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_avg_price_cmd_lastIdx       : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_avg_price_cmd_ctrl          : out std_logic_vector(L_AVG_PRICE_BUS_ADDR_WIDTH - 1 downto 0);
      l_avg_price_cmd_tag           : out std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_avg_disc_cmd_valid          : out std_logic;
      l_avg_disc_cmd_ready          : in std_logic;
      l_avg_disc_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_avg_disc_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_avg_disc_cmd_ctrl           : out std_logic_vector(L_AVG_DISC_BUS_ADDR_WIDTH - 1 downto 0);
      l_avg_disc_cmd_tag            : out std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_count_order_cmd_valid       : out std_logic;
      l_count_order_cmd_ready       : in std_logic;
      l_count_order_cmd_firstIdx    : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_count_order_cmd_lastIdx     : out std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_count_order_cmd_ctrl        : out std_logic_vector(L_COUNT_ORDER_BUS_ADDR_WIDTH - 1 downto 0);
      l_count_order_cmd_tag         : out std_logic_vector(TAG_WIDTH - 1 downto 0)

    );
  end component;

  component PriceSummary_l is
    generic (
      INDEX_WIDTH                         : integer := 32;
      TAG_WIDTH                           : integer := 1;
      L_QUANTITY_BUS_ADDR_WIDTH           : integer := 64;
      L_QUANTITY_BUS_DATA_WIDTH           : integer := 512;
      L_QUANTITY_BUS_LEN_WIDTH            : integer := 8;
      L_QUANTITY_BUS_BURST_STEP_LEN       : integer := 1;
      L_QUANTITY_BUS_BURST_MAX_LEN        : integer := 16;
      L_EXTENDEDPRICE_BUS_ADDR_WIDTH      : integer := 64;
      L_EXTENDEDPRICE_BUS_DATA_WIDTH      : integer := 512;
      L_EXTENDEDPRICE_BUS_LEN_WIDTH       : integer := 8;
      L_EXTENDEDPRICE_BUS_BURST_STEP_LEN  : integer := 1;
      L_EXTENDEDPRICE_BUS_BURST_MAX_LEN   : integer := 16;
      L_DISCOUNT_BUS_ADDR_WIDTH           : integer := 64;
      L_DISCOUNT_BUS_DATA_WIDTH           : integer := 512;
      L_DISCOUNT_BUS_LEN_WIDTH            : integer := 8;
      L_DISCOUNT_BUS_BURST_STEP_LEN       : integer := 1;
      L_DISCOUNT_BUS_BURST_MAX_LEN        : integer := 16;
      L_TAX_BUS_ADDR_WIDTH                : integer := 64;
      L_TAX_BUS_DATA_WIDTH                : integer := 512;
      L_TAX_BUS_LEN_WIDTH                 : integer := 8;
      L_TAX_BUS_BURST_STEP_LEN            : integer := 1;
      L_TAX_BUS_BURST_MAX_LEN             : integer := 16;
      L_RETURNFLAG_BUS_ADDR_WIDTH         : integer := 64;
      L_RETURNFLAG_BUS_DATA_WIDTH         : integer := 512;
      L_RETURNFLAG_BUS_LEN_WIDTH          : integer := 8;
      L_RETURNFLAG_BUS_BURST_STEP_LEN     : integer := 1;
      L_RETURNFLAG_BUS_BURST_MAX_LEN      : integer := 16;
      L_LINESTATUS_BUS_ADDR_WIDTH         : integer := 64;
      L_LINESTATUS_BUS_DATA_WIDTH         : integer := 512;
      L_LINESTATUS_BUS_LEN_WIDTH          : integer := 8;
      L_LINESTATUS_BUS_BURST_STEP_LEN     : integer := 1;
      L_LINESTATUS_BUS_BURST_MAX_LEN      : integer := 16;
      L_SHIPDATE_BUS_ADDR_WIDTH           : integer := 64;
      L_SHIPDATE_BUS_DATA_WIDTH           : integer := 512;
      L_SHIPDATE_BUS_LEN_WIDTH            : integer := 8;
      L_SHIPDATE_BUS_BURST_STEP_LEN       : integer := 1;
      L_SHIPDATE_BUS_BURST_MAX_LEN        : integer := 16;
      L_RETURNFLAG_O_BUS_ADDR_WIDTH       : integer := 64;
      L_RETURNFLAG_O_BUS_DATA_WIDTH       : integer := 512;
      L_RETURNFLAG_O_BUS_LEN_WIDTH        : integer := 8;
      L_RETURNFLAG_O_BUS_BURST_STEP_LEN   : integer := 1;
      L_RETURNFLAG_O_BUS_BURST_MAX_LEN    : integer := 16;
      L_LINESTATUS_O_BUS_ADDR_WIDTH       : integer := 64;
      L_LINESTATUS_O_BUS_DATA_WIDTH       : integer := 512;
      L_LINESTATUS_O_BUS_LEN_WIDTH        : integer := 8;
      L_LINESTATUS_O_BUS_BURST_STEP_LEN   : integer := 1;
      L_LINESTATUS_O_BUS_BURST_MAX_LEN    : integer := 16;
      L_SUM_QTY_BUS_ADDR_WIDTH            : integer := 64;
      L_SUM_QTY_BUS_DATA_WIDTH            : integer := 512;
      L_SUM_QTY_BUS_LEN_WIDTH             : integer := 8;
      L_SUM_QTY_BUS_BURST_STEP_LEN        : integer := 1;
      L_SUM_QTY_BUS_BURST_MAX_LEN         : integer := 16;
      L_SUM_BASE_PRICE_BUS_ADDR_WIDTH     : integer := 64;
      L_SUM_BASE_PRICE_BUS_DATA_WIDTH     : integer := 512;
      L_SUM_BASE_PRICE_BUS_LEN_WIDTH      : integer := 8;
      L_SUM_BASE_PRICE_BUS_BURST_STEP_LEN : integer := 1;
      L_SUM_BASE_PRICE_BUS_BURST_MAX_LEN  : integer := 16;
      L_SUM_DISC_PRICE_BUS_ADDR_WIDTH     : integer := 64;
      L_SUM_DISC_PRICE_BUS_DATA_WIDTH     : integer := 512;
      L_SUM_DISC_PRICE_BUS_LEN_WIDTH      : integer := 8;
      L_SUM_DISC_PRICE_BUS_BURST_STEP_LEN : integer := 1;
      L_SUM_DISC_PRICE_BUS_BURST_MAX_LEN  : integer := 16;
      L_SUM_CHARGE_BUS_ADDR_WIDTH         : integer := 64;
      L_SUM_CHARGE_BUS_DATA_WIDTH         : integer := 512;
      L_SUM_CHARGE_BUS_LEN_WIDTH          : integer := 8;
      L_SUM_CHARGE_BUS_BURST_STEP_LEN     : integer := 1;
      L_SUM_CHARGE_BUS_BURST_MAX_LEN      : integer := 16;
      L_AVG_QTY_BUS_ADDR_WIDTH            : integer := 64;
      L_AVG_QTY_BUS_DATA_WIDTH            : integer := 512;
      L_AVG_QTY_BUS_LEN_WIDTH             : integer := 8;
      L_AVG_QTY_BUS_BURST_STEP_LEN        : integer := 1;
      L_AVG_QTY_BUS_BURST_MAX_LEN         : integer := 16;
      L_AVG_PRICE_BUS_ADDR_WIDTH          : integer := 64;
      L_AVG_PRICE_BUS_DATA_WIDTH          : integer := 512;
      L_AVG_PRICE_BUS_LEN_WIDTH           : integer := 8;
      L_AVG_PRICE_BUS_BURST_STEP_LEN      : integer := 1;
      L_AVG_PRICE_BUS_BURST_MAX_LEN       : integer := 16;
      L_AVG_DISC_BUS_ADDR_WIDTH           : integer := 64;
      L_AVG_DISC_BUS_DATA_WIDTH           : integer := 512;
      L_AVG_DISC_BUS_LEN_WIDTH            : integer := 8;
      L_AVG_DISC_BUS_BURST_STEP_LEN       : integer := 1;
      L_AVG_DISC_BUS_BURST_MAX_LEN        : integer := 16;
      L_COUNT_ORDER_BUS_ADDR_WIDTH        : integer := 64;
      L_COUNT_ORDER_BUS_DATA_WIDTH        : integer := 512;
      L_COUNT_ORDER_BUS_LEN_WIDTH         : integer := 8;
      L_COUNT_ORDER_BUS_BURST_STEP_LEN    : integer := 1;
      L_COUNT_ORDER_BUS_BURST_MAX_LEN     : integer := 16
    );
    port (
      bcd_clk                          : in std_logic;
      bcd_reset                        : in std_logic;
      kcd_clk                          : in std_logic;
      kcd_reset                        : in std_logic;
      l_quantity_valid                 : out std_logic;
      l_quantity_ready                 : in std_logic;
      l_quantity_dvalid                : out std_logic;
      l_quantity_last                  : out std_logic;
      l_quantity                       : out std_logic_vector(63 downto 0);
      l_quantity_bus_rreq_valid        : out std_logic;
      l_quantity_bus_rreq_ready        : in std_logic;
      l_quantity_bus_rreq_addr         : out std_logic_vector(L_QUANTITY_BUS_ADDR_WIDTH - 1 downto 0);
      l_quantity_bus_rreq_len          : out std_logic_vector(L_QUANTITY_BUS_LEN_WIDTH - 1 downto 0);
      l_quantity_bus_rdat_valid        : in std_logic;
      l_quantity_bus_rdat_ready        : out std_logic;
      l_quantity_bus_rdat_data         : in std_logic_vector(L_QUANTITY_BUS_DATA_WIDTH - 1 downto 0);
      l_quantity_bus_rdat_last         : in std_logic;
      l_quantity_cmd_valid             : in std_logic;
      l_quantity_cmd_ready             : out std_logic;
      l_quantity_cmd_firstIdx          : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_quantity_cmd_lastIdx           : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_quantity_cmd_ctrl              : in std_logic_vector(L_QUANTITY_BUS_ADDR_WIDTH - 1 downto 0);
      l_quantity_cmd_tag               : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_quantity_unl_valid             : out std_logic;
      l_quantity_unl_ready             : in std_logic;
      l_quantity_unl_tag               : out std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_extendedprice_valid            : out std_logic;
      l_extendedprice_ready            : in std_logic;
      l_extendedprice_dvalid           : out std_logic;
      l_extendedprice_last             : out std_logic;
      l_extendedprice                  : out std_logic_vector(63 downto 0);
      l_extendedprice_bus_rreq_valid   : out std_logic;
      l_extendedprice_bus_rreq_ready   : in std_logic;
      l_extendedprice_bus_rreq_addr    : out std_logic_vector(L_EXTENDEDPRICE_BUS_ADDR_WIDTH - 1 downto 0);
      l_extendedprice_bus_rreq_len     : out std_logic_vector(L_EXTENDEDPRICE_BUS_LEN_WIDTH - 1 downto 0);
      l_extendedprice_bus_rdat_valid   : in std_logic;
      l_extendedprice_bus_rdat_ready   : out std_logic;
      l_extendedprice_bus_rdat_data    : in std_logic_vector(L_EXTENDEDPRICE_BUS_DATA_WIDTH - 1 downto 0);
      l_extendedprice_bus_rdat_last    : in std_logic;
      l_extendedprice_cmd_valid        : in std_logic;
      l_extendedprice_cmd_ready        : out std_logic;
      l_extendedprice_cmd_firstIdx     : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_extendedprice_cmd_lastIdx      : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_extendedprice_cmd_ctrl         : in std_logic_vector(L_EXTENDEDPRICE_BUS_ADDR_WIDTH - 1 downto 0);
      l_extendedprice_cmd_tag          : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_extendedprice_unl_valid        : out std_logic;
      l_extendedprice_unl_ready        : in std_logic;
      l_extendedprice_unl_tag          : out std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_discount_valid                 : out std_logic;
      l_discount_ready                 : in std_logic;
      l_discount_dvalid                : out std_logic;
      l_discount_last                  : out std_logic;
      l_discount                       : out std_logic_vector(63 downto 0);
      l_discount_bus_rreq_valid        : out std_logic;
      l_discount_bus_rreq_ready        : in std_logic;
      l_discount_bus_rreq_addr         : out std_logic_vector(L_DISCOUNT_BUS_ADDR_WIDTH - 1 downto 0);
      l_discount_bus_rreq_len          : out std_logic_vector(L_DISCOUNT_BUS_LEN_WIDTH - 1 downto 0);
      l_discount_bus_rdat_valid        : in std_logic;
      l_discount_bus_rdat_ready        : out std_logic;
      l_discount_bus_rdat_data         : in std_logic_vector(L_DISCOUNT_BUS_DATA_WIDTH - 1 downto 0);
      l_discount_bus_rdat_last         : in std_logic;
      l_discount_cmd_valid             : in std_logic;
      l_discount_cmd_ready             : out std_logic;
      l_discount_cmd_firstIdx          : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_discount_cmd_lastIdx           : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_discount_cmd_ctrl              : in std_logic_vector(L_DISCOUNT_BUS_ADDR_WIDTH - 1 downto 0);
      l_discount_cmd_tag               : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_discount_unl_valid             : out std_logic;
      l_discount_unl_ready             : in std_logic;
      l_discount_unl_tag               : out std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_tax_valid                      : out std_logic;
      l_tax_ready                      : in std_logic;
      l_tax_dvalid                     : out std_logic;
      l_tax_last                       : out std_logic;
      l_tax                            : out std_logic_vector(63 downto 0);
      l_tax_bus_rreq_valid             : out std_logic;
      l_tax_bus_rreq_ready             : in std_logic;
      l_tax_bus_rreq_addr              : out std_logic_vector(L_TAX_BUS_ADDR_WIDTH - 1 downto 0);
      l_tax_bus_rreq_len               : out std_logic_vector(L_TAX_BUS_LEN_WIDTH - 1 downto 0);
      l_tax_bus_rdat_valid             : in std_logic;
      l_tax_bus_rdat_ready             : out std_logic;
      l_tax_bus_rdat_data              : in std_logic_vector(L_TAX_BUS_DATA_WIDTH - 1 downto 0);
      l_tax_bus_rdat_last              : in std_logic;
      l_tax_cmd_valid                  : in std_logic;
      l_tax_cmd_ready                  : out std_logic;
      l_tax_cmd_firstIdx               : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_tax_cmd_lastIdx                : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_tax_cmd_ctrl                   : in std_logic_vector(L_TAX_BUS_ADDR_WIDTH - 1 downto 0);
      l_tax_cmd_tag                    : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_tax_unl_valid                  : out std_logic;
      l_tax_unl_ready                  : in std_logic;
      l_tax_unl_tag                    : out std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_returnflag_valid               : out std_logic;
      l_returnflag_ready               : in std_logic;
      l_returnflag_dvalid              : out std_logic;
      l_returnflag_last                : out std_logic;
      l_returnflag_length              : out std_logic_vector(31 downto 0);
      l_returnflag_count               : out std_logic_vector(0 downto 0);
      l_returnflag_chars_valid         : out std_logic;
      l_returnflag_chars_ready         : in std_logic;
      l_returnflag_chars_dvalid        : out std_logic;
      l_returnflag_chars_last          : out std_logic;
      l_returnflag_chars               : out std_logic_vector(7 downto 0);
      l_returnflag_chars_count         : out std_logic_vector(0 downto 0);
      l_returnflag_bus_rreq_valid      : out std_logic;
      l_returnflag_bus_rreq_ready      : in std_logic;
      l_returnflag_bus_rreq_addr       : out std_logic_vector(L_RETURNFLAG_BUS_ADDR_WIDTH - 1 downto 0);
      l_returnflag_bus_rreq_len        : out std_logic_vector(L_RETURNFLAG_BUS_LEN_WIDTH - 1 downto 0);
      l_returnflag_bus_rdat_valid      : in std_logic;
      l_returnflag_bus_rdat_ready      : out std_logic;
      l_returnflag_bus_rdat_data       : in std_logic_vector(L_RETURNFLAG_BUS_DATA_WIDTH - 1 downto 0);
      l_returnflag_bus_rdat_last       : in std_logic;
      l_returnflag_cmd_valid           : in std_logic;
      l_returnflag_cmd_ready           : out std_logic;
      l_returnflag_cmd_firstIdx        : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_returnflag_cmd_lastIdx         : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_returnflag_cmd_ctrl            : in std_logic_vector(L_RETURNFLAG_BUS_ADDR_WIDTH * 2 - 1 downto 0);
      l_returnflag_cmd_tag             : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_returnflag_unl_valid           : out std_logic;
      l_returnflag_unl_ready           : in std_logic;
      l_returnflag_unl_tag             : out std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_linestatus_valid               : out std_logic;
      l_linestatus_ready               : in std_logic;
      l_linestatus_dvalid              : out std_logic;
      l_linestatus_last                : out std_logic;
      l_linestatus_length              : out std_logic_vector(31 downto 0);
      l_linestatus_count               : out std_logic_vector(0 downto 0);
      l_linestatus_chars_valid         : out std_logic;
      l_linestatus_chars_ready         : in std_logic;
      l_linestatus_chars_dvalid        : out std_logic;
      l_linestatus_chars_last          : out std_logic;
      l_linestatus_chars               : out std_logic_vector(7 downto 0);
      l_linestatus_chars_count         : out std_logic_vector(0 downto 0);
      l_linestatus_bus_rreq_valid      : out std_logic;
      l_linestatus_bus_rreq_ready      : in std_logic;
      l_linestatus_bus_rreq_addr       : out std_logic_vector(L_LINESTATUS_BUS_ADDR_WIDTH - 1 downto 0);
      l_linestatus_bus_rreq_len        : out std_logic_vector(L_LINESTATUS_BUS_LEN_WIDTH - 1 downto 0);
      l_linestatus_bus_rdat_valid      : in std_logic;
      l_linestatus_bus_rdat_ready      : out std_logic;
      l_linestatus_bus_rdat_data       : in std_logic_vector(L_LINESTATUS_BUS_DATA_WIDTH - 1 downto 0);
      l_linestatus_bus_rdat_last       : in std_logic;
      l_linestatus_cmd_valid           : in std_logic;
      l_linestatus_cmd_ready           : out std_logic;
      l_linestatus_cmd_firstIdx        : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_linestatus_cmd_lastIdx         : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_linestatus_cmd_ctrl            : in std_logic_vector(L_LINESTATUS_BUS_ADDR_WIDTH * 2 - 1 downto 0);
      l_linestatus_cmd_tag             : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_linestatus_unl_valid           : out std_logic;
      l_linestatus_unl_ready           : in std_logic;
      l_linestatus_unl_tag             : out std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_shipdate_valid                 : out std_logic;
      l_shipdate_ready                 : in std_logic;
      l_shipdate_dvalid                : out std_logic;
      l_shipdate_last                  : out std_logic;
      l_shipdate                       : out std_logic_vector(31 downto 0);
      l_shipdate_bus_rreq_valid        : out std_logic;
      l_shipdate_bus_rreq_ready        : in std_logic;
      l_shipdate_bus_rreq_addr         : out std_logic_vector(L_SHIPDATE_BUS_ADDR_WIDTH - 1 downto 0);
      l_shipdate_bus_rreq_len          : out std_logic_vector(L_SHIPDATE_BUS_LEN_WIDTH - 1 downto 0);
      l_shipdate_bus_rdat_valid        : in std_logic;
      l_shipdate_bus_rdat_ready        : out std_logic;
      l_shipdate_bus_rdat_data         : in std_logic_vector(L_SHIPDATE_BUS_DATA_WIDTH - 1 downto 0);
      l_shipdate_bus_rdat_last         : in std_logic;
      l_shipdate_cmd_valid             : in std_logic;
      l_shipdate_cmd_ready             : out std_logic;
      l_shipdate_cmd_firstIdx          : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_shipdate_cmd_lastIdx           : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_shipdate_cmd_ctrl              : in std_logic_vector(L_SHIPDATE_BUS_ADDR_WIDTH - 1 downto 0);
      l_shipdate_cmd_tag               : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_shipdate_unl_valid             : out std_logic;
      l_shipdate_unl_ready             : in std_logic;
      l_shipdate_unl_tag               : out std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_returnflag_o_valid             : in std_logic;
      l_returnflag_o_ready             : out std_logic;
      l_returnflag_o_dvalid            : in std_logic;
      l_returnflag_o_last              : in std_logic;
      l_returnflag_o_length            : in std_logic_vector(31 downto 0);
      l_returnflag_o_count             : in std_logic_vector(0 downto 0);
      l_returnflag_o_chars_valid       : in std_logic;
      l_returnflag_o_chars_ready       : out std_logic;
      l_returnflag_o_chars_dvalid      : in std_logic;
      l_returnflag_o_chars_last        : in std_logic;
      l_returnflag_o_chars             : in std_logic_vector(7 downto 0);
      l_returnflag_o_chars_count       : in std_logic_vector(0 downto 0);
      l_returnflag_o_bus_wreq_valid    : out std_logic;
      l_returnflag_o_bus_wreq_ready    : in std_logic;
      l_returnflag_o_bus_wreq_addr     : out std_logic_vector(L_RETURNFLAG_O_BUS_ADDR_WIDTH - 1 downto 0);
      l_returnflag_o_bus_wreq_len      : out std_logic_vector(L_RETURNFLAG_O_BUS_LEN_WIDTH - 1 downto 0);
      l_returnflag_o_bus_wdat_valid    : out std_logic;
      l_returnflag_o_bus_wdat_ready    : in std_logic;
      l_returnflag_o_bus_wdat_data     : out std_logic_vector(L_RETURNFLAG_O_BUS_DATA_WIDTH - 1 downto 0);
      l_returnflag_o_bus_wdat_strobe   : out std_logic_vector(L_RETURNFLAG_O_BUS_DATA_WIDTH/8 - 1 downto 0);
      l_returnflag_o_bus_wdat_last     : out std_logic;
      l_returnflag_o_cmd_valid         : in std_logic;
      l_returnflag_o_cmd_ready         : out std_logic;
      l_returnflag_o_cmd_firstIdx      : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_returnflag_o_cmd_lastIdx       : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_returnflag_o_cmd_ctrl          : in std_logic_vector(L_RETURNFLAG_O_BUS_ADDR_WIDTH * 2 - 1 downto 0);
      l_returnflag_o_cmd_tag           : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_returnflag_o_unl_valid         : out std_logic;
      l_returnflag_o_unl_ready         : in std_logic;
      l_returnflag_o_unl_tag           : out std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_linestatus_o_valid             : in std_logic;
      l_linestatus_o_ready             : out std_logic;
      l_linestatus_o_dvalid            : in std_logic;
      l_linestatus_o_last              : in std_logic;
      l_linestatus_o_length            : in std_logic_vector(31 downto 0);
      l_linestatus_o_count             : in std_logic_vector(0 downto 0);
      l_linestatus_o_chars_valid       : in std_logic;
      l_linestatus_o_chars_ready       : out std_logic;
      l_linestatus_o_chars_dvalid      : in std_logic;
      l_linestatus_o_chars_last        : in std_logic;
      l_linestatus_o_chars             : in std_logic_vector(7 downto 0);
      l_linestatus_o_chars_count       : in std_logic_vector(0 downto 0);
      l_linestatus_o_bus_wreq_valid    : out std_logic;
      l_linestatus_o_bus_wreq_ready    : in std_logic;
      l_linestatus_o_bus_wreq_addr     : out std_logic_vector(L_LINESTATUS_O_BUS_ADDR_WIDTH - 1 downto 0);
      l_linestatus_o_bus_wreq_len      : out std_logic_vector(L_LINESTATUS_O_BUS_LEN_WIDTH - 1 downto 0);
      l_linestatus_o_bus_wdat_valid    : out std_logic;
      l_linestatus_o_bus_wdat_ready    : in std_logic;
      l_linestatus_o_bus_wdat_data     : out std_logic_vector(L_LINESTATUS_O_BUS_DATA_WIDTH - 1 downto 0);
      l_linestatus_o_bus_wdat_strobe   : out std_logic_vector(L_LINESTATUS_O_BUS_DATA_WIDTH/8 - 1 downto 0);
      l_linestatus_o_bus_wdat_last     : out std_logic;
      l_linestatus_o_cmd_valid         : in std_logic;
      l_linestatus_o_cmd_ready         : out std_logic;
      l_linestatus_o_cmd_firstIdx      : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_linestatus_o_cmd_lastIdx       : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_linestatus_o_cmd_ctrl          : in std_logic_vector(L_LINESTATUS_O_BUS_ADDR_WIDTH * 2 - 1 downto 0);
      l_linestatus_o_cmd_tag           : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_linestatus_o_unl_valid         : out std_logic;
      l_linestatus_o_unl_ready         : in std_logic;
      l_linestatus_o_unl_tag           : out std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_sum_qty_valid                  : in std_logic;
      l_sum_qty_ready                  : out std_logic;
      l_sum_qty_dvalid                 : in std_logic;
      l_sum_qty_last                   : in std_logic;
      l_sum_qty                        : in std_logic_vector(63 downto 0);
      l_sum_qty_bus_wreq_valid         : out std_logic;
      l_sum_qty_bus_wreq_ready         : in std_logic;
      l_sum_qty_bus_wreq_addr          : out std_logic_vector(L_SUM_QTY_BUS_ADDR_WIDTH - 1 downto 0);
      l_sum_qty_bus_wreq_len           : out std_logic_vector(L_SUM_QTY_BUS_LEN_WIDTH - 1 downto 0);
      l_sum_qty_bus_wdat_valid         : out std_logic;
      l_sum_qty_bus_wdat_ready         : in std_logic;
      l_sum_qty_bus_wdat_data          : out std_logic_vector(L_SUM_QTY_BUS_DATA_WIDTH - 1 downto 0);
      l_sum_qty_bus_wdat_strobe        : out std_logic_vector(L_SUM_QTY_BUS_DATA_WIDTH/8 - 1 downto 0);
      l_sum_qty_bus_wdat_last          : out std_logic;
      l_sum_qty_cmd_valid              : in std_logic;
      l_sum_qty_cmd_ready              : out std_logic;
      l_sum_qty_cmd_firstIdx           : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_sum_qty_cmd_lastIdx            : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_sum_qty_cmd_ctrl               : in std_logic_vector(L_SUM_QTY_BUS_ADDR_WIDTH - 1 downto 0);
      l_sum_qty_cmd_tag                : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_sum_qty_unl_valid              : out std_logic;
      l_sum_qty_unl_ready              : in std_logic;
      l_sum_qty_unl_tag                : out std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_sum_base_price_valid           : in std_logic;
      l_sum_base_price_ready           : out std_logic;
      l_sum_base_price_dvalid          : in std_logic;
      l_sum_base_price_last            : in std_logic;
      l_sum_base_price                 : in std_logic_vector(63 downto 0);
      l_sum_base_price_bus_wreq_valid  : out std_logic;
      l_sum_base_price_bus_wreq_ready  : in std_logic;
      l_sum_base_price_bus_wreq_addr   : out std_logic_vector(L_SUM_BASE_PRICE_BUS_ADDR_WIDTH - 1 downto 0);
      l_sum_base_price_bus_wreq_len    : out std_logic_vector(L_SUM_BASE_PRICE_BUS_LEN_WIDTH - 1 downto 0);
      l_sum_base_price_bus_wdat_valid  : out std_logic;
      l_sum_base_price_bus_wdat_ready  : in std_logic;
      l_sum_base_price_bus_wdat_data   : out std_logic_vector(L_SUM_BASE_PRICE_BUS_DATA_WIDTH - 1 downto 0);
      l_sum_base_price_bus_wdat_strobe : out std_logic_vector(L_SUM_BASE_PRICE_BUS_DATA_WIDTH/8 - 1 downto 0);
      l_sum_base_price_bus_wdat_last   : out std_logic;
      l_sum_base_price_cmd_valid       : in std_logic;
      l_sum_base_price_cmd_ready       : out std_logic;
      l_sum_base_price_cmd_firstIdx    : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_sum_base_price_cmd_lastIdx     : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_sum_base_price_cmd_ctrl        : in std_logic_vector(L_SUM_BASE_PRICE_BUS_ADDR_WIDTH - 1 downto 0);
      l_sum_base_price_cmd_tag         : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_sum_base_price_unl_valid       : out std_logic;
      l_sum_base_price_unl_ready       : in std_logic;
      l_sum_base_price_unl_tag         : out std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_sum_disc_price_valid           : in std_logic;
      l_sum_disc_price_ready           : out std_logic;
      l_sum_disc_price_dvalid          : in std_logic;
      l_sum_disc_price_last            : in std_logic;
      l_sum_disc_price                 : in std_logic_vector(63 downto 0);
      l_sum_disc_price_bus_wreq_valid  : out std_logic;
      l_sum_disc_price_bus_wreq_ready  : in std_logic;
      l_sum_disc_price_bus_wreq_addr   : out std_logic_vector(L_SUM_DISC_PRICE_BUS_ADDR_WIDTH - 1 downto 0);
      l_sum_disc_price_bus_wreq_len    : out std_logic_vector(L_SUM_DISC_PRICE_BUS_LEN_WIDTH - 1 downto 0);
      l_sum_disc_price_bus_wdat_valid  : out std_logic;
      l_sum_disc_price_bus_wdat_ready  : in std_logic;
      l_sum_disc_price_bus_wdat_data   : out std_logic_vector(L_SUM_DISC_PRICE_BUS_DATA_WIDTH - 1 downto 0);
      l_sum_disc_price_bus_wdat_strobe : out std_logic_vector(L_SUM_DISC_PRICE_BUS_DATA_WIDTH/8 - 1 downto 0);
      l_sum_disc_price_bus_wdat_last   : out std_logic;
      l_sum_disc_price_cmd_valid       : in std_logic;
      l_sum_disc_price_cmd_ready       : out std_logic;
      l_sum_disc_price_cmd_firstIdx    : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_sum_disc_price_cmd_lastIdx     : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_sum_disc_price_cmd_ctrl        : in std_logic_vector(L_SUM_DISC_PRICE_BUS_ADDR_WIDTH - 1 downto 0);
      l_sum_disc_price_cmd_tag         : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_sum_disc_price_unl_valid       : out std_logic;
      l_sum_disc_price_unl_ready       : in std_logic;
      l_sum_disc_price_unl_tag         : out std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_sum_charge_valid               : in std_logic;
      l_sum_charge_ready               : out std_logic;
      l_sum_charge_dvalid              : in std_logic;
      l_sum_charge_last                : in std_logic;
      l_sum_charge                     : in std_logic_vector(63 downto 0);
      l_sum_charge_bus_wreq_valid      : out std_logic;
      l_sum_charge_bus_wreq_ready      : in std_logic;
      l_sum_charge_bus_wreq_addr       : out std_logic_vector(L_SUM_CHARGE_BUS_ADDR_WIDTH - 1 downto 0);
      l_sum_charge_bus_wreq_len        : out std_logic_vector(L_SUM_CHARGE_BUS_LEN_WIDTH - 1 downto 0);
      l_sum_charge_bus_wdat_valid      : out std_logic;
      l_sum_charge_bus_wdat_ready      : in std_logic;
      l_sum_charge_bus_wdat_data       : out std_logic_vector(L_SUM_CHARGE_BUS_DATA_WIDTH - 1 downto 0);
      l_sum_charge_bus_wdat_strobe     : out std_logic_vector(L_SUM_CHARGE_BUS_DATA_WIDTH/8 - 1 downto 0);
      l_sum_charge_bus_wdat_last       : out std_logic;
      l_sum_charge_cmd_valid           : in std_logic;
      l_sum_charge_cmd_ready           : out std_logic;
      l_sum_charge_cmd_firstIdx        : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_sum_charge_cmd_lastIdx         : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_sum_charge_cmd_ctrl            : in std_logic_vector(L_SUM_CHARGE_BUS_ADDR_WIDTH - 1 downto 0);
      l_sum_charge_cmd_tag             : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_sum_charge_unl_valid           : out std_logic;
      l_sum_charge_unl_ready           : in std_logic;
      l_sum_charge_unl_tag             : out std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_avg_qty_valid                  : in std_logic;
      l_avg_qty_ready                  : out std_logic;
      l_avg_qty_dvalid                 : in std_logic;
      l_avg_qty_last                   : in std_logic;
      l_avg_qty                        : in std_logic_vector(63 downto 0);
      l_avg_qty_bus_wreq_valid         : out std_logic;
      l_avg_qty_bus_wreq_ready         : in std_logic;
      l_avg_qty_bus_wreq_addr          : out std_logic_vector(L_AVG_QTY_BUS_ADDR_WIDTH - 1 downto 0);
      l_avg_qty_bus_wreq_len           : out std_logic_vector(L_AVG_QTY_BUS_LEN_WIDTH - 1 downto 0);
      l_avg_qty_bus_wdat_valid         : out std_logic;
      l_avg_qty_bus_wdat_ready         : in std_logic;
      l_avg_qty_bus_wdat_data          : out std_logic_vector(L_AVG_QTY_BUS_DATA_WIDTH - 1 downto 0);
      l_avg_qty_bus_wdat_strobe        : out std_logic_vector(L_AVG_QTY_BUS_DATA_WIDTH/8 - 1 downto 0);
      l_avg_qty_bus_wdat_last          : out std_logic;
      l_avg_qty_cmd_valid              : in std_logic;
      l_avg_qty_cmd_ready              : out std_logic;
      l_avg_qty_cmd_firstIdx           : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_avg_qty_cmd_lastIdx            : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_avg_qty_cmd_ctrl               : in std_logic_vector(L_AVG_QTY_BUS_ADDR_WIDTH - 1 downto 0);
      l_avg_qty_cmd_tag                : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_avg_qty_unl_valid              : out std_logic;
      l_avg_qty_unl_ready              : in std_logic;
      l_avg_qty_unl_tag                : out std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_avg_price_valid                : in std_logic;
      l_avg_price_ready                : out std_logic;
      l_avg_price_dvalid               : in std_logic;
      l_avg_price_last                 : in std_logic;
      l_avg_price                      : in std_logic_vector(63 downto 0);
      l_avg_price_bus_wreq_valid       : out std_logic;
      l_avg_price_bus_wreq_ready       : in std_logic;
      l_avg_price_bus_wreq_addr        : out std_logic_vector(L_AVG_PRICE_BUS_ADDR_WIDTH - 1 downto 0);
      l_avg_price_bus_wreq_len         : out std_logic_vector(L_AVG_PRICE_BUS_LEN_WIDTH - 1 downto 0);
      l_avg_price_bus_wdat_valid       : out std_logic;
      l_avg_price_bus_wdat_ready       : in std_logic;
      l_avg_price_bus_wdat_data        : out std_logic_vector(L_AVG_PRICE_BUS_DATA_WIDTH - 1 downto 0);
      l_avg_price_bus_wdat_strobe      : out std_logic_vector(L_AVG_PRICE_BUS_DATA_WIDTH/8 - 1 downto 0);
      l_avg_price_bus_wdat_last        : out std_logic;
      l_avg_price_cmd_valid            : in std_logic;
      l_avg_price_cmd_ready            : out std_logic;
      l_avg_price_cmd_firstIdx         : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_avg_price_cmd_lastIdx          : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_avg_price_cmd_ctrl             : in std_logic_vector(L_AVG_PRICE_BUS_ADDR_WIDTH - 1 downto 0);
      l_avg_price_cmd_tag              : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_avg_price_unl_valid            : out std_logic;
      l_avg_price_unl_ready            : in std_logic;
      l_avg_price_unl_tag              : out std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_avg_disc_valid                 : in std_logic;
      l_avg_disc_ready                 : out std_logic;
      l_avg_disc_dvalid                : in std_logic;
      l_avg_disc_last                  : in std_logic;
      l_avg_disc                       : in std_logic_vector(63 downto 0);
      l_avg_disc_bus_wreq_valid        : out std_logic;
      l_avg_disc_bus_wreq_ready        : in std_logic;
      l_avg_disc_bus_wreq_addr         : out std_logic_vector(L_AVG_DISC_BUS_ADDR_WIDTH - 1 downto 0);
      l_avg_disc_bus_wreq_len          : out std_logic_vector(L_AVG_DISC_BUS_LEN_WIDTH - 1 downto 0);
      l_avg_disc_bus_wdat_valid        : out std_logic;
      l_avg_disc_bus_wdat_ready        : in std_logic;
      l_avg_disc_bus_wdat_data         : out std_logic_vector(L_AVG_DISC_BUS_DATA_WIDTH - 1 downto 0);
      l_avg_disc_bus_wdat_strobe       : out std_logic_vector(L_AVG_DISC_BUS_DATA_WIDTH/8 - 1 downto 0);
      l_avg_disc_bus_wdat_last         : out std_logic;
      l_avg_disc_cmd_valid             : in std_logic;
      l_avg_disc_cmd_ready             : out std_logic;
      l_avg_disc_cmd_firstIdx          : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_avg_disc_cmd_lastIdx           : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_avg_disc_cmd_ctrl              : in std_logic_vector(L_AVG_DISC_BUS_ADDR_WIDTH - 1 downto 0);
      l_avg_disc_cmd_tag               : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_avg_disc_unl_valid             : out std_logic;
      l_avg_disc_unl_ready             : in std_logic;
      l_avg_disc_unl_tag               : out std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_count_order_valid              : in std_logic;
      l_count_order_ready              : out std_logic;
      l_count_order_dvalid             : in std_logic;
      l_count_order_last               : in std_logic;
      l_count_order                    : in std_logic_vector(63 downto 0);
      l_count_order_bus_wreq_valid     : out std_logic;
      l_count_order_bus_wreq_ready     : in std_logic;
      l_count_order_bus_wreq_addr      : out std_logic_vector(L_COUNT_ORDER_BUS_ADDR_WIDTH - 1 downto 0);
      l_count_order_bus_wreq_len       : out std_logic_vector(L_COUNT_ORDER_BUS_LEN_WIDTH - 1 downto 0);
      l_count_order_bus_wdat_valid     : out std_logic;
      l_count_order_bus_wdat_ready     : in std_logic;
      l_count_order_bus_wdat_data      : out std_logic_vector(L_COUNT_ORDER_BUS_DATA_WIDTH - 1 downto 0);
      l_count_order_bus_wdat_strobe    : out std_logic_vector(L_COUNT_ORDER_BUS_DATA_WIDTH/8 - 1 downto 0);
      l_count_order_bus_wdat_last      : out std_logic;
      l_count_order_cmd_valid          : in std_logic;
      l_count_order_cmd_ready          : out std_logic;
      l_count_order_cmd_firstIdx       : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_count_order_cmd_lastIdx        : in std_logic_vector(INDEX_WIDTH - 1 downto 0);
      l_count_order_cmd_ctrl           : in std_logic_vector(L_COUNT_ORDER_BUS_ADDR_WIDTH - 1 downto 0);
      l_count_order_cmd_tag            : in std_logic_vector(TAG_WIDTH - 1 downto 0);
      l_count_order_unl_valid          : out std_logic;
      l_count_order_unl_ready          : in std_logic;
      l_count_order_unl_tag            : out std_logic_vector(TAG_WIDTH - 1 downto 0)
    );
  end component;

  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_valid          : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_ready          : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_dvalid         : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_last           : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_length         : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_count          : std_logic_vector(0 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_valid    : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_ready    : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_dvalid   : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_last     : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars          : std_logic_vector(7 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_count    : std_logic_vector(0 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_valid          : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_ready          : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_dvalid         : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_last           : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_length         : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_count          : std_logic_vector(0 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_valid    : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_ready    : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_dvalid   : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_last     : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars          : std_logic_vector(7 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_count    : std_logic_vector(0 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_sum_qty_valid               : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_qty_ready               : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_qty_dvalid              : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_qty_last                : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_qty                     : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_sum_base_price_valid        : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_base_price_ready        : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_base_price_dvalid       : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_base_price_last         : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_base_price              : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_valid        : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_ready        : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_dvalid       : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_last         : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_disc_price              : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_sum_charge_valid            : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_charge_ready            : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_charge_dvalid           : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_charge_last             : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_charge                  : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_avg_qty_valid               : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_qty_ready               : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_qty_dvalid              : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_qty_last                : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_qty                     : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_avg_price_valid             : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_price_ready             : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_price_dvalid            : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_price_last              : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_price                   : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_avg_disc_valid              : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_disc_ready              : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_disc_dvalid             : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_disc_last               : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_disc                    : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_count_order_valid           : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_count_order_ready           : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_count_order_dvalid          : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_count_order_last            : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_count_order                 : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_unl_valid      : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_unl_ready      : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_unl_tag        : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_unl_valid      : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_unl_ready      : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_unl_tag        : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_sum_qty_unl_valid           : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_qty_unl_ready           : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_qty_unl_tag             : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_sum_base_price_unl_valid    : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_base_price_unl_ready    : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_base_price_unl_tag      : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_unl_valid    : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_unl_ready    : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_unl_tag      : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_sum_charge_unl_valid        : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_charge_unl_ready        : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_charge_unl_tag          : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_avg_qty_unl_valid           : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_qty_unl_ready           : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_qty_unl_tag             : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_avg_price_unl_valid         : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_price_unl_ready         : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_price_unl_tag           : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_avg_disc_unl_valid          : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_disc_unl_ready          : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_disc_unl_tag            : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_count_order_unl_valid       : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_count_order_unl_ready       : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_count_order_unl_tag         : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_valid      : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_ready      : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_firstIdx   : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_lastIdx    : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_ctrl       : std_logic_vector(BUS_ADDR_WIDTH * 2 - 1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_tag        : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_valid      : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_ready      : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_firstIdx   : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_lastIdx    : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_ctrl       : std_logic_vector(BUS_ADDR_WIDTH * 2 - 1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_tag        : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_valid           : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_ready           : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_firstIdx        : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_lastIdx         : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_ctrl            : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_tag             : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_valid    : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_ready    : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_firstIdx : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_lastIdx  : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_ctrl     : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_tag      : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_valid    : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_ready    : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_firstIdx : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_lastIdx  : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_ctrl     : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_tag      : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_valid        : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_ready        : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_firstIdx     : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_lastIdx      : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_ctrl         : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_tag          : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_valid           : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_ready           : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_firstIdx        : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_lastIdx         : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_ctrl            : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_tag             : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_valid         : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_ready         : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_ctrl          : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_tag           : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_valid          : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_ready          : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_ctrl           : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_tag            : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_valid       : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_ready       : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_firstIdx    : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_lastIdx     : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_ctrl        : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_tag         : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_l_inst_l_returnflag_o_valid                : std_logic;
  signal PriceSummaryWriter_l_inst_l_returnflag_o_ready                : std_logic;
  signal PriceSummaryWriter_l_inst_l_returnflag_o_dvalid               : std_logic;
  signal PriceSummaryWriter_l_inst_l_returnflag_o_last                 : std_logic;
  signal PriceSummaryWriter_l_inst_l_returnflag_o_length               : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_l_inst_l_returnflag_o_count                : std_logic_vector(0 downto 0);
  signal PriceSummaryWriter_l_inst_l_returnflag_o_chars_valid          : std_logic;
  signal PriceSummaryWriter_l_inst_l_returnflag_o_chars_ready          : std_logic;
  signal PriceSummaryWriter_l_inst_l_returnflag_o_chars_dvalid         : std_logic;
  signal PriceSummaryWriter_l_inst_l_returnflag_o_chars_last           : std_logic;
  signal PriceSummaryWriter_l_inst_l_returnflag_o_chars                : std_logic_vector(7 downto 0);
  signal PriceSummaryWriter_l_inst_l_returnflag_o_chars_count          : std_logic_vector(0 downto 0);

  signal PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_valid       : std_logic;
  signal PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_ready       : std_logic;
  signal PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_addr        : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_len         : std_logic_vector(BUS_LEN_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_valid       : std_logic;
  signal PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_ready       : std_logic;
  signal PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_data        : std_logic_vector(BUS_DATA_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_strobe      : std_logic_vector(BUS_DATA_WIDTH/8 - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_last        : std_logic;

  signal PriceSummaryWriter_l_inst_l_returnflag_o_cmd_valid            : std_logic;
  signal PriceSummaryWriter_l_inst_l_returnflag_o_cmd_ready            : std_logic;
  signal PriceSummaryWriter_l_inst_l_returnflag_o_cmd_firstIdx         : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_returnflag_o_cmd_lastIdx          : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_returnflag_o_cmd_ctrl             : std_logic_vector(BUS_ADDR_WIDTH * 2 - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_returnflag_o_cmd_tag              : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_l_inst_l_returnflag_o_unl_valid            : std_logic;
  signal PriceSummaryWriter_l_inst_l_returnflag_o_unl_ready            : std_logic;
  signal PriceSummaryWriter_l_inst_l_returnflag_o_unl_tag              : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_l_inst_l_linestatus_o_valid                : std_logic;
  signal PriceSummaryWriter_l_inst_l_linestatus_o_ready                : std_logic;
  signal PriceSummaryWriter_l_inst_l_linestatus_o_dvalid               : std_logic;
  signal PriceSummaryWriter_l_inst_l_linestatus_o_last                 : std_logic;
  signal PriceSummaryWriter_l_inst_l_linestatus_o_length               : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_l_inst_l_linestatus_o_count                : std_logic_vector(0 downto 0);
  signal PriceSummaryWriter_l_inst_l_linestatus_o_chars_valid          : std_logic;
  signal PriceSummaryWriter_l_inst_l_linestatus_o_chars_ready          : std_logic;
  signal PriceSummaryWriter_l_inst_l_linestatus_o_chars_dvalid         : std_logic;
  signal PriceSummaryWriter_l_inst_l_linestatus_o_chars_last           : std_logic;
  signal PriceSummaryWriter_l_inst_l_linestatus_o_chars                : std_logic_vector(7 downto 0);
  signal PriceSummaryWriter_l_inst_l_linestatus_o_chars_count          : std_logic_vector(0 downto 0);

  signal PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_valid       : std_logic;
  signal PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_ready       : std_logic;
  signal PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_addr        : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_len         : std_logic_vector(BUS_LEN_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_valid       : std_logic;
  signal PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_ready       : std_logic;
  signal PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_data        : std_logic_vector(BUS_DATA_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_strobe      : std_logic_vector(BUS_DATA_WIDTH/8 - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_last        : std_logic;

  signal PriceSummaryWriter_l_inst_l_linestatus_o_cmd_valid            : std_logic;
  signal PriceSummaryWriter_l_inst_l_linestatus_o_cmd_ready            : std_logic;
  signal PriceSummaryWriter_l_inst_l_linestatus_o_cmd_firstIdx         : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_linestatus_o_cmd_lastIdx          : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_linestatus_o_cmd_ctrl             : std_logic_vector(BUS_ADDR_WIDTH * 2 - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_linestatus_o_cmd_tag              : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_l_inst_l_linestatus_o_unl_valid            : std_logic;
  signal PriceSummaryWriter_l_inst_l_linestatus_o_unl_ready            : std_logic;
  signal PriceSummaryWriter_l_inst_l_linestatus_o_unl_tag              : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_l_inst_l_sum_qty_valid                     : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_qty_ready                     : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_qty_dvalid                    : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_qty_last                      : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_qty                           : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_valid            : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_ready            : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_addr             : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_len              : std_logic_vector(BUS_LEN_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_valid            : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_ready            : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_data             : std_logic_vector(BUS_DATA_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_strobe           : std_logic_vector(BUS_DATA_WIDTH/8 - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_last             : std_logic;

  signal PriceSummaryWriter_l_inst_l_sum_qty_cmd_valid                 : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_qty_cmd_ready                 : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_qty_cmd_firstIdx              : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_qty_cmd_lastIdx               : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_qty_cmd_ctrl                  : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_qty_cmd_tag                   : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_l_inst_l_sum_qty_unl_valid                 : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_qty_unl_ready                 : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_qty_unl_tag                   : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_l_inst_l_sum_base_price_valid              : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_base_price_ready              : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_base_price_dvalid             : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_base_price_last               : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_base_price                    : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_valid     : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_ready     : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_addr      : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_len       : std_logic_vector(BUS_LEN_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_valid     : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_ready     : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_data      : std_logic_vector(BUS_DATA_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_strobe    : std_logic_vector(BUS_DATA_WIDTH/8 - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_last      : std_logic;

  signal PriceSummaryWriter_l_inst_l_sum_base_price_cmd_valid          : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_base_price_cmd_ready          : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_base_price_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_base_price_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_base_price_cmd_ctrl           : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_base_price_cmd_tag            : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_l_inst_l_sum_base_price_unl_valid          : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_base_price_unl_ready          : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_base_price_unl_tag            : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_l_inst_l_sum_disc_price_valid              : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_ready              : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_dvalid             : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_last               : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_disc_price                    : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_valid     : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_ready     : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_addr      : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_len       : std_logic_vector(BUS_LEN_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_valid     : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_ready     : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_data      : std_logic_vector(BUS_DATA_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_strobe    : std_logic_vector(BUS_DATA_WIDTH/8 - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_last      : std_logic;

  signal PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_valid          : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_ready          : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_ctrl           : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_tag            : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_l_inst_l_sum_disc_price_unl_valid          : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_unl_ready          : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_unl_tag            : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_l_inst_l_sum_charge_valid                  : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_charge_ready                  : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_charge_dvalid                 : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_charge_last                   : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_charge                        : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_valid         : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_ready         : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_addr          : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_len           : std_logic_vector(BUS_LEN_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_valid         : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_ready         : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_data          : std_logic_vector(BUS_DATA_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_strobe        : std_logic_vector(BUS_DATA_WIDTH/8 - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_last          : std_logic;

  signal PriceSummaryWriter_l_inst_l_sum_charge_cmd_valid              : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_charge_cmd_ready              : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_charge_cmd_firstIdx           : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_charge_cmd_lastIdx            : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_charge_cmd_ctrl               : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_charge_cmd_tag                : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_l_inst_l_sum_charge_unl_valid              : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_charge_unl_ready              : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_charge_unl_tag                : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_l_inst_l_avg_qty_valid                     : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_qty_ready                     : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_qty_dvalid                    : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_qty_last                      : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_qty                           : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_valid            : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_ready            : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_addr             : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_len              : std_logic_vector(BUS_LEN_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_valid            : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_ready            : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_data             : std_logic_vector(BUS_DATA_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_strobe           : std_logic_vector(BUS_DATA_WIDTH/8 - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_last             : std_logic;

  signal PriceSummaryWriter_l_inst_l_avg_qty_cmd_valid                 : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_qty_cmd_ready                 : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_qty_cmd_firstIdx              : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_qty_cmd_lastIdx               : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_qty_cmd_ctrl                  : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_qty_cmd_tag                   : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_l_inst_l_avg_qty_unl_valid                 : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_qty_unl_ready                 : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_qty_unl_tag                   : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_l_inst_l_avg_price_valid                   : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_price_ready                   : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_price_dvalid                  : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_price_last                    : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_price                         : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_valid          : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_ready          : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_addr           : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_len            : std_logic_vector(BUS_LEN_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_valid          : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_ready          : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_data           : std_logic_vector(BUS_DATA_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_strobe         : std_logic_vector(BUS_DATA_WIDTH/8 - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_last           : std_logic;

  signal PriceSummaryWriter_l_inst_l_avg_price_cmd_valid               : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_price_cmd_ready               : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_price_cmd_firstIdx            : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_price_cmd_lastIdx             : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_price_cmd_ctrl                : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_price_cmd_tag                 : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_l_inst_l_avg_price_unl_valid               : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_price_unl_ready               : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_price_unl_tag                 : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_l_inst_l_avg_disc_valid                    : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_disc_ready                    : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_disc_dvalid                   : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_disc_last                     : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_disc                          : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_valid           : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_ready           : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_addr            : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_len             : std_logic_vector(BUS_LEN_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_valid           : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_ready           : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_data            : std_logic_vector(BUS_DATA_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_strobe          : std_logic_vector(BUS_DATA_WIDTH/8 - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_last            : std_logic;

  signal PriceSummaryWriter_l_inst_l_avg_disc_cmd_valid                : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_disc_cmd_ready                : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_disc_cmd_firstIdx             : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_disc_cmd_lastIdx              : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_disc_cmd_ctrl                 : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_disc_cmd_tag                  : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_l_inst_l_avg_disc_unl_valid                : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_disc_unl_ready                : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_disc_unl_tag                  : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_l_inst_l_count_order_valid                 : std_logic;
  signal PriceSummaryWriter_l_inst_l_count_order_ready                 : std_logic;
  signal PriceSummaryWriter_l_inst_l_count_order_dvalid                : std_logic;
  signal PriceSummaryWriter_l_inst_l_count_order_last                  : std_logic;
  signal PriceSummaryWriter_l_inst_l_count_order                       : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_l_inst_l_count_order_bus_wreq_valid        : std_logic;
  signal PriceSummaryWriter_l_inst_l_count_order_bus_wreq_ready        : std_logic;
  signal PriceSummaryWriter_l_inst_l_count_order_bus_wreq_addr         : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_count_order_bus_wreq_len          : std_logic_vector(BUS_LEN_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_count_order_bus_wdat_valid        : std_logic;
  signal PriceSummaryWriter_l_inst_l_count_order_bus_wdat_ready        : std_logic;
  signal PriceSummaryWriter_l_inst_l_count_order_bus_wdat_data         : std_logic_vector(BUS_DATA_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_count_order_bus_wdat_strobe       : std_logic_vector(BUS_DATA_WIDTH/8 - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_count_order_bus_wdat_last         : std_logic;

  signal PriceSummaryWriter_l_inst_l_count_order_cmd_valid             : std_logic;
  signal PriceSummaryWriter_l_inst_l_count_order_cmd_ready             : std_logic;
  signal PriceSummaryWriter_l_inst_l_count_order_cmd_firstIdx          : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_count_order_cmd_lastIdx           : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_count_order_cmd_ctrl              : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummaryWriter_l_inst_l_count_order_cmd_tag               : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummaryWriter_l_inst_l_count_order_unl_valid             : std_logic;
  signal PriceSummaryWriter_l_inst_l_count_order_unl_ready             : std_logic;
  signal PriceSummaryWriter_l_inst_l_count_order_unl_tag               : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummary_Nucleus_inst_mmio_awvalid                        : std_logic;
  signal PriceSummary_Nucleus_inst_mmio_awready                        : std_logic;
  signal PriceSummary_Nucleus_inst_mmio_awaddr                         : std_logic_vector(31 downto 0);
  signal PriceSummary_Nucleus_inst_mmio_wvalid                         : std_logic;
  signal PriceSummary_Nucleus_inst_mmio_wready                         : std_logic;
  signal PriceSummary_Nucleus_inst_mmio_wdata                          : std_logic_vector(31 downto 0);
  signal PriceSummary_Nucleus_inst_mmio_wstrb                          : std_logic_vector(3 downto 0);
  signal PriceSummary_Nucleus_inst_mmio_bvalid                         : std_logic;
  signal PriceSummary_Nucleus_inst_mmio_bready                         : std_logic;
  signal PriceSummary_Nucleus_inst_mmio_bresp                          : std_logic_vector(1 downto 0);
  signal PriceSummary_Nucleus_inst_mmio_arvalid                        : std_logic;
  signal PriceSummary_Nucleus_inst_mmio_arready                        : std_logic;
  signal PriceSummary_Nucleus_inst_mmio_araddr                         : std_logic_vector(31 downto 0);
  signal PriceSummary_Nucleus_inst_mmio_rvalid                         : std_logic;
  signal PriceSummary_Nucleus_inst_mmio_rready                         : std_logic;
  signal PriceSummary_Nucleus_inst_mmio_rdata                          : std_logic_vector(31 downto 0);
  signal PriceSummary_Nucleus_inst_mmio_rresp                          : std_logic_vector(1 downto 0);

  signal PriceSummary_Nucleus_inst_l_quantity_valid                    : std_logic;
  signal PriceSummary_Nucleus_inst_l_quantity_ready                    : std_logic;
  signal PriceSummary_Nucleus_inst_l_quantity_dvalid                   : std_logic;
  signal PriceSummary_Nucleus_inst_l_quantity_last                     : std_logic;
  signal PriceSummary_Nucleus_inst_l_quantity                          : std_logic_vector(63 downto 0);

  signal PriceSummary_Nucleus_inst_l_extendedprice_valid               : std_logic;
  signal PriceSummary_Nucleus_inst_l_extendedprice_ready               : std_logic;
  signal PriceSummary_Nucleus_inst_l_extendedprice_dvalid              : std_logic;
  signal PriceSummary_Nucleus_inst_l_extendedprice_last                : std_logic;
  signal PriceSummary_Nucleus_inst_l_extendedprice                     : std_logic_vector(63 downto 0);

  signal PriceSummary_Nucleus_inst_l_discount_valid                    : std_logic;
  signal PriceSummary_Nucleus_inst_l_discount_ready                    : std_logic;
  signal PriceSummary_Nucleus_inst_l_discount_dvalid                   : std_logic;
  signal PriceSummary_Nucleus_inst_l_discount_last                     : std_logic;
  signal PriceSummary_Nucleus_inst_l_discount                          : std_logic_vector(63 downto 0);

  signal PriceSummary_Nucleus_inst_l_tax_valid                         : std_logic;
  signal PriceSummary_Nucleus_inst_l_tax_ready                         : std_logic;
  signal PriceSummary_Nucleus_inst_l_tax_dvalid                        : std_logic;
  signal PriceSummary_Nucleus_inst_l_tax_last                          : std_logic;
  signal PriceSummary_Nucleus_inst_l_tax                               : std_logic_vector(63 downto 0);

  signal PriceSummary_Nucleus_inst_l_returnflag_valid                  : std_logic;
  signal PriceSummary_Nucleus_inst_l_returnflag_ready                  : std_logic;
  signal PriceSummary_Nucleus_inst_l_returnflag_dvalid                 : std_logic;
  signal PriceSummary_Nucleus_inst_l_returnflag_last                   : std_logic;
  signal PriceSummary_Nucleus_inst_l_returnflag_length                 : std_logic_vector(31 downto 0);
  signal PriceSummary_Nucleus_inst_l_returnflag_count                  : std_logic_vector(0 downto 0);
  signal PriceSummary_Nucleus_inst_l_returnflag_chars_valid            : std_logic;
  signal PriceSummary_Nucleus_inst_l_returnflag_chars_ready            : std_logic;
  signal PriceSummary_Nucleus_inst_l_returnflag_chars_dvalid           : std_logic;
  signal PriceSummary_Nucleus_inst_l_returnflag_chars_last             : std_logic;
  signal PriceSummary_Nucleus_inst_l_returnflag_chars                  : std_logic_vector(7 downto 0);
  signal PriceSummary_Nucleus_inst_l_returnflag_chars_count            : std_logic_vector(0 downto 0);

  signal PriceSummary_Nucleus_inst_l_linestatus_valid                  : std_logic;
  signal PriceSummary_Nucleus_inst_l_linestatus_ready                  : std_logic;
  signal PriceSummary_Nucleus_inst_l_linestatus_dvalid                 : std_logic;
  signal PriceSummary_Nucleus_inst_l_linestatus_last                   : std_logic;
  signal PriceSummary_Nucleus_inst_l_linestatus_length                 : std_logic_vector(31 downto 0);
  signal PriceSummary_Nucleus_inst_l_linestatus_count                  : std_logic_vector(0 downto 0);
  signal PriceSummary_Nucleus_inst_l_linestatus_chars_valid            : std_logic;
  signal PriceSummary_Nucleus_inst_l_linestatus_chars_ready            : std_logic;
  signal PriceSummary_Nucleus_inst_l_linestatus_chars_dvalid           : std_logic;
  signal PriceSummary_Nucleus_inst_l_linestatus_chars_last             : std_logic;
  signal PriceSummary_Nucleus_inst_l_linestatus_chars                  : std_logic_vector(7 downto 0);
  signal PriceSummary_Nucleus_inst_l_linestatus_chars_count            : std_logic_vector(0 downto 0);

  signal PriceSummary_Nucleus_inst_l_shipdate_valid                    : std_logic;
  signal PriceSummary_Nucleus_inst_l_shipdate_ready                    : std_logic;
  signal PriceSummary_Nucleus_inst_l_shipdate_dvalid                   : std_logic;
  signal PriceSummary_Nucleus_inst_l_shipdate_last                     : std_logic;
  signal PriceSummary_Nucleus_inst_l_shipdate                          : std_logic_vector(31 downto 0);

  signal PriceSummary_Nucleus_inst_l_quantity_unl_valid                : std_logic;
  signal PriceSummary_Nucleus_inst_l_quantity_unl_ready                : std_logic;
  signal PriceSummary_Nucleus_inst_l_quantity_unl_tag                  : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummary_Nucleus_inst_l_extendedprice_unl_valid           : std_logic;
  signal PriceSummary_Nucleus_inst_l_extendedprice_unl_ready           : std_logic;
  signal PriceSummary_Nucleus_inst_l_extendedprice_unl_tag             : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummary_Nucleus_inst_l_discount_unl_valid                : std_logic;
  signal PriceSummary_Nucleus_inst_l_discount_unl_ready                : std_logic;
  signal PriceSummary_Nucleus_inst_l_discount_unl_tag                  : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummary_Nucleus_inst_l_tax_unl_valid                     : std_logic;
  signal PriceSummary_Nucleus_inst_l_tax_unl_ready                     : std_logic;
  signal PriceSummary_Nucleus_inst_l_tax_unl_tag                       : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummary_Nucleus_inst_l_returnflag_unl_valid              : std_logic;
  signal PriceSummary_Nucleus_inst_l_returnflag_unl_ready              : std_logic;
  signal PriceSummary_Nucleus_inst_l_returnflag_unl_tag                : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummary_Nucleus_inst_l_linestatus_unl_valid              : std_logic;
  signal PriceSummary_Nucleus_inst_l_linestatus_unl_ready              : std_logic;
  signal PriceSummary_Nucleus_inst_l_linestatus_unl_tag                : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummary_Nucleus_inst_l_shipdate_unl_valid                : std_logic;
  signal PriceSummary_Nucleus_inst_l_shipdate_unl_ready                : std_logic;
  signal PriceSummary_Nucleus_inst_l_shipdate_unl_tag                  : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummary_Nucleus_inst_l_quantity_cmd_valid                : std_logic;
  signal PriceSummary_Nucleus_inst_l_quantity_cmd_ready                : std_logic;
  signal PriceSummary_Nucleus_inst_l_quantity_cmd_firstIdx             : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummary_Nucleus_inst_l_quantity_cmd_lastIdx              : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummary_Nucleus_inst_l_quantity_cmd_ctrl                 : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummary_Nucleus_inst_l_quantity_cmd_tag                  : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummary_Nucleus_inst_l_extendedprice_cmd_valid           : std_logic;
  signal PriceSummary_Nucleus_inst_l_extendedprice_cmd_ready           : std_logic;
  signal PriceSummary_Nucleus_inst_l_extendedprice_cmd_firstIdx        : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummary_Nucleus_inst_l_extendedprice_cmd_lastIdx         : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummary_Nucleus_inst_l_extendedprice_cmd_ctrl            : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummary_Nucleus_inst_l_extendedprice_cmd_tag             : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummary_Nucleus_inst_l_discount_cmd_valid                : std_logic;
  signal PriceSummary_Nucleus_inst_l_discount_cmd_ready                : std_logic;
  signal PriceSummary_Nucleus_inst_l_discount_cmd_firstIdx             : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummary_Nucleus_inst_l_discount_cmd_lastIdx              : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummary_Nucleus_inst_l_discount_cmd_ctrl                 : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummary_Nucleus_inst_l_discount_cmd_tag                  : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummary_Nucleus_inst_l_tax_cmd_valid                     : std_logic;
  signal PriceSummary_Nucleus_inst_l_tax_cmd_ready                     : std_logic;
  signal PriceSummary_Nucleus_inst_l_tax_cmd_firstIdx                  : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummary_Nucleus_inst_l_tax_cmd_lastIdx                   : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummary_Nucleus_inst_l_tax_cmd_ctrl                      : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummary_Nucleus_inst_l_tax_cmd_tag                       : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummary_Nucleus_inst_l_returnflag_cmd_valid              : std_logic;
  signal PriceSummary_Nucleus_inst_l_returnflag_cmd_ready              : std_logic;
  signal PriceSummary_Nucleus_inst_l_returnflag_cmd_firstIdx           : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummary_Nucleus_inst_l_returnflag_cmd_lastIdx            : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummary_Nucleus_inst_l_returnflag_cmd_ctrl               : std_logic_vector(BUS_ADDR_WIDTH * 2 - 1 downto 0);
  signal PriceSummary_Nucleus_inst_l_returnflag_cmd_tag                : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummary_Nucleus_inst_l_linestatus_cmd_valid              : std_logic;
  signal PriceSummary_Nucleus_inst_l_linestatus_cmd_ready              : std_logic;
  signal PriceSummary_Nucleus_inst_l_linestatus_cmd_firstIdx           : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummary_Nucleus_inst_l_linestatus_cmd_lastIdx            : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummary_Nucleus_inst_l_linestatus_cmd_ctrl               : std_logic_vector(BUS_ADDR_WIDTH * 2 - 1 downto 0);
  signal PriceSummary_Nucleus_inst_l_linestatus_cmd_tag                : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummary_Nucleus_inst_l_shipdate_cmd_valid                : std_logic;
  signal PriceSummary_Nucleus_inst_l_shipdate_cmd_ready                : std_logic;
  signal PriceSummary_Nucleus_inst_l_shipdate_cmd_firstIdx             : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummary_Nucleus_inst_l_shipdate_cmd_lastIdx              : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummary_Nucleus_inst_l_shipdate_cmd_ctrl                 : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummary_Nucleus_inst_l_shipdate_cmd_tag                  : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummary_l_inst_l_quantity_valid                          : std_logic;
  signal PriceSummary_l_inst_l_quantity_ready                          : std_logic;
  signal PriceSummary_l_inst_l_quantity_dvalid                         : std_logic;
  signal PriceSummary_l_inst_l_quantity_last                           : std_logic;
  signal PriceSummary_l_inst_l_quantity                                : std_logic_vector(63 downto 0);

  signal PriceSummary_l_inst_l_quantity_bus_rreq_valid                 : std_logic;
  signal PriceSummary_l_inst_l_quantity_bus_rreq_ready                 : std_logic;
  signal PriceSummary_l_inst_l_quantity_bus_rreq_addr                  : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_quantity_bus_rreq_len                   : std_logic_vector(BUS_LEN_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_quantity_bus_rdat_valid                 : std_logic;
  signal PriceSummary_l_inst_l_quantity_bus_rdat_ready                 : std_logic;
  signal PriceSummary_l_inst_l_quantity_bus_rdat_data                  : std_logic_vector(BUS_DATA_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_quantity_bus_rdat_last                  : std_logic;

  signal PriceSummary_l_inst_l_quantity_cmd_valid                      : std_logic;
  signal PriceSummary_l_inst_l_quantity_cmd_ready                      : std_logic;
  signal PriceSummary_l_inst_l_quantity_cmd_firstIdx                   : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_quantity_cmd_lastIdx                    : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_quantity_cmd_ctrl                       : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_quantity_cmd_tag                        : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummary_l_inst_l_quantity_unl_valid                      : std_logic;
  signal PriceSummary_l_inst_l_quantity_unl_ready                      : std_logic;
  signal PriceSummary_l_inst_l_quantity_unl_tag                        : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummary_l_inst_l_extendedprice_valid                     : std_logic;
  signal PriceSummary_l_inst_l_extendedprice_ready                     : std_logic;
  signal PriceSummary_l_inst_l_extendedprice_dvalid                    : std_logic;
  signal PriceSummary_l_inst_l_extendedprice_last                      : std_logic;
  signal PriceSummary_l_inst_l_extendedprice                           : std_logic_vector(63 downto 0);

  signal PriceSummary_l_inst_l_extendedprice_bus_rreq_valid            : std_logic;
  signal PriceSummary_l_inst_l_extendedprice_bus_rreq_ready            : std_logic;
  signal PriceSummary_l_inst_l_extendedprice_bus_rreq_addr             : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_extendedprice_bus_rreq_len              : std_logic_vector(BUS_LEN_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_extendedprice_bus_rdat_valid            : std_logic;
  signal PriceSummary_l_inst_l_extendedprice_bus_rdat_ready            : std_logic;
  signal PriceSummary_l_inst_l_extendedprice_bus_rdat_data             : std_logic_vector(BUS_DATA_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_extendedprice_bus_rdat_last             : std_logic;

  signal PriceSummary_l_inst_l_extendedprice_cmd_valid                 : std_logic;
  signal PriceSummary_l_inst_l_extendedprice_cmd_ready                 : std_logic;
  signal PriceSummary_l_inst_l_extendedprice_cmd_firstIdx              : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_extendedprice_cmd_lastIdx               : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_extendedprice_cmd_ctrl                  : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_extendedprice_cmd_tag                   : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummary_l_inst_l_extendedprice_unl_valid                 : std_logic;
  signal PriceSummary_l_inst_l_extendedprice_unl_ready                 : std_logic;
  signal PriceSummary_l_inst_l_extendedprice_unl_tag                   : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummary_l_inst_l_discount_valid                          : std_logic;
  signal PriceSummary_l_inst_l_discount_ready                          : std_logic;
  signal PriceSummary_l_inst_l_discount_dvalid                         : std_logic;
  signal PriceSummary_l_inst_l_discount_last                           : std_logic;
  signal PriceSummary_l_inst_l_discount                                : std_logic_vector(63 downto 0);

  signal PriceSummary_l_inst_l_discount_bus_rreq_valid                 : std_logic;
  signal PriceSummary_l_inst_l_discount_bus_rreq_ready                 : std_logic;
  signal PriceSummary_l_inst_l_discount_bus_rreq_addr                  : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_discount_bus_rreq_len                   : std_logic_vector(BUS_LEN_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_discount_bus_rdat_valid                 : std_logic;
  signal PriceSummary_l_inst_l_discount_bus_rdat_ready                 : std_logic;
  signal PriceSummary_l_inst_l_discount_bus_rdat_data                  : std_logic_vector(BUS_DATA_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_discount_bus_rdat_last                  : std_logic;

  signal PriceSummary_l_inst_l_discount_cmd_valid                      : std_logic;
  signal PriceSummary_l_inst_l_discount_cmd_ready                      : std_logic;
  signal PriceSummary_l_inst_l_discount_cmd_firstIdx                   : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_discount_cmd_lastIdx                    : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_discount_cmd_ctrl                       : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_discount_cmd_tag                        : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummary_l_inst_l_discount_unl_valid                      : std_logic;
  signal PriceSummary_l_inst_l_discount_unl_ready                      : std_logic;
  signal PriceSummary_l_inst_l_discount_unl_tag                        : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummary_l_inst_l_tax_valid                               : std_logic;
  signal PriceSummary_l_inst_l_tax_ready                               : std_logic;
  signal PriceSummary_l_inst_l_tax_dvalid                              : std_logic;
  signal PriceSummary_l_inst_l_tax_last                                : std_logic;
  signal PriceSummary_l_inst_l_tax                                     : std_logic_vector(63 downto 0);

  signal PriceSummary_l_inst_l_tax_bus_rreq_valid                      : std_logic;
  signal PriceSummary_l_inst_l_tax_bus_rreq_ready                      : std_logic;
  signal PriceSummary_l_inst_l_tax_bus_rreq_addr                       : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_tax_bus_rreq_len                        : std_logic_vector(BUS_LEN_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_tax_bus_rdat_valid                      : std_logic;
  signal PriceSummary_l_inst_l_tax_bus_rdat_ready                      : std_logic;
  signal PriceSummary_l_inst_l_tax_bus_rdat_data                       : std_logic_vector(BUS_DATA_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_tax_bus_rdat_last                       : std_logic;

  signal PriceSummary_l_inst_l_tax_cmd_valid                           : std_logic;
  signal PriceSummary_l_inst_l_tax_cmd_ready                           : std_logic;
  signal PriceSummary_l_inst_l_tax_cmd_firstIdx                        : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_tax_cmd_lastIdx                         : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_tax_cmd_ctrl                            : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_tax_cmd_tag                             : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummary_l_inst_l_tax_unl_valid                           : std_logic;
  signal PriceSummary_l_inst_l_tax_unl_ready                           : std_logic;
  signal PriceSummary_l_inst_l_tax_unl_tag                             : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummary_l_inst_l_returnflag_valid                        : std_logic;
  signal PriceSummary_l_inst_l_returnflag_ready                        : std_logic;
  signal PriceSummary_l_inst_l_returnflag_dvalid                       : std_logic;
  signal PriceSummary_l_inst_l_returnflag_last                         : std_logic;
  signal PriceSummary_l_inst_l_returnflag_length                       : std_logic_vector(31 downto 0);
  signal PriceSummary_l_inst_l_returnflag_count                        : std_logic_vector(0 downto 0);
  signal PriceSummary_l_inst_l_returnflag_chars_valid                  : std_logic;
  signal PriceSummary_l_inst_l_returnflag_chars_ready                  : std_logic;
  signal PriceSummary_l_inst_l_returnflag_chars_dvalid                 : std_logic;
  signal PriceSummary_l_inst_l_returnflag_chars_last                   : std_logic;
  signal PriceSummary_l_inst_l_returnflag_chars                        : std_logic_vector(7 downto 0);
  signal PriceSummary_l_inst_l_returnflag_chars_count                  : std_logic_vector(0 downto 0);

  signal PriceSummary_l_inst_l_returnflag_bus_rreq_valid               : std_logic;
  signal PriceSummary_l_inst_l_returnflag_bus_rreq_ready               : std_logic;
  signal PriceSummary_l_inst_l_returnflag_bus_rreq_addr                : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_returnflag_bus_rreq_len                 : std_logic_vector(BUS_LEN_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_returnflag_bus_rdat_valid               : std_logic;
  signal PriceSummary_l_inst_l_returnflag_bus_rdat_ready               : std_logic;
  signal PriceSummary_l_inst_l_returnflag_bus_rdat_data                : std_logic_vector(BUS_DATA_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_returnflag_bus_rdat_last                : std_logic;

  signal PriceSummary_l_inst_l_returnflag_cmd_valid                    : std_logic;
  signal PriceSummary_l_inst_l_returnflag_cmd_ready                    : std_logic;
  signal PriceSummary_l_inst_l_returnflag_cmd_firstIdx                 : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_returnflag_cmd_lastIdx                  : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_returnflag_cmd_ctrl                     : std_logic_vector(BUS_ADDR_WIDTH * 2 - 1 downto 0);
  signal PriceSummary_l_inst_l_returnflag_cmd_tag                      : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummary_l_inst_l_returnflag_unl_valid                    : std_logic;
  signal PriceSummary_l_inst_l_returnflag_unl_ready                    : std_logic;
  signal PriceSummary_l_inst_l_returnflag_unl_tag                      : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummary_l_inst_l_linestatus_valid                        : std_logic;
  signal PriceSummary_l_inst_l_linestatus_ready                        : std_logic;
  signal PriceSummary_l_inst_l_linestatus_dvalid                       : std_logic;
  signal PriceSummary_l_inst_l_linestatus_last                         : std_logic;
  signal PriceSummary_l_inst_l_linestatus_length                       : std_logic_vector(31 downto 0);
  signal PriceSummary_l_inst_l_linestatus_count                        : std_logic_vector(0 downto 0);
  signal PriceSummary_l_inst_l_linestatus_chars_valid                  : std_logic;
  signal PriceSummary_l_inst_l_linestatus_chars_ready                  : std_logic;
  signal PriceSummary_l_inst_l_linestatus_chars_dvalid                 : std_logic;
  signal PriceSummary_l_inst_l_linestatus_chars_last                   : std_logic;
  signal PriceSummary_l_inst_l_linestatus_chars                        : std_logic_vector(7 downto 0);
  signal PriceSummary_l_inst_l_linestatus_chars_count                  : std_logic_vector(0 downto 0);

  signal PriceSummary_l_inst_l_linestatus_bus_rreq_valid               : std_logic;
  signal PriceSummary_l_inst_l_linestatus_bus_rreq_ready               : std_logic;
  signal PriceSummary_l_inst_l_linestatus_bus_rreq_addr                : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_linestatus_bus_rreq_len                 : std_logic_vector(BUS_LEN_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_linestatus_bus_rdat_valid               : std_logic;
  signal PriceSummary_l_inst_l_linestatus_bus_rdat_ready               : std_logic;
  signal PriceSummary_l_inst_l_linestatus_bus_rdat_data                : std_logic_vector(BUS_DATA_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_linestatus_bus_rdat_last                : std_logic;

  signal PriceSummary_l_inst_l_linestatus_cmd_valid                    : std_logic;
  signal PriceSummary_l_inst_l_linestatus_cmd_ready                    : std_logic;
  signal PriceSummary_l_inst_l_linestatus_cmd_firstIdx                 : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_linestatus_cmd_lastIdx                  : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_linestatus_cmd_ctrl                     : std_logic_vector(BUS_ADDR_WIDTH * 2 - 1 downto 0);
  signal PriceSummary_l_inst_l_linestatus_cmd_tag                      : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummary_l_inst_l_linestatus_unl_valid                    : std_logic;
  signal PriceSummary_l_inst_l_linestatus_unl_ready                    : std_logic;
  signal PriceSummary_l_inst_l_linestatus_unl_tag                      : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummary_l_inst_l_shipdate_valid                          : std_logic;
  signal PriceSummary_l_inst_l_shipdate_ready                          : std_logic;
  signal PriceSummary_l_inst_l_shipdate_dvalid                         : std_logic;
  signal PriceSummary_l_inst_l_shipdate_last                           : std_logic;
  signal PriceSummary_l_inst_l_shipdate                                : std_logic_vector(31 downto 0);

  signal PriceSummary_l_inst_l_shipdate_bus_rreq_valid                 : std_logic;
  signal PriceSummary_l_inst_l_shipdate_bus_rreq_ready                 : std_logic;
  signal PriceSummary_l_inst_l_shipdate_bus_rreq_addr                  : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_shipdate_bus_rreq_len                   : std_logic_vector(BUS_LEN_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_shipdate_bus_rdat_valid                 : std_logic;
  signal PriceSummary_l_inst_l_shipdate_bus_rdat_ready                 : std_logic;
  signal PriceSummary_l_inst_l_shipdate_bus_rdat_data                  : std_logic_vector(BUS_DATA_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_shipdate_bus_rdat_last                  : std_logic;

  signal PriceSummary_l_inst_l_shipdate_cmd_valid                      : std_logic;
  signal PriceSummary_l_inst_l_shipdate_cmd_ready                      : std_logic;
  signal PriceSummary_l_inst_l_shipdate_cmd_firstIdx                   : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_shipdate_cmd_lastIdx                    : std_logic_vector(INDEX_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_shipdate_cmd_ctrl                       : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal PriceSummary_l_inst_l_shipdate_cmd_tag                        : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal PriceSummary_l_inst_l_shipdate_unl_valid                      : std_logic;
  signal PriceSummary_l_inst_l_shipdate_unl_ready                      : std_logic;
  signal PriceSummary_l_inst_l_shipdate_unl_tag                        : std_logic_vector(TAG_WIDTH - 1 downto 0);

  signal RDAW64DW512LW8BS1BM16_inst_mst_rreq_valid                     : std_logic;
  signal RDAW64DW512LW8BS1BM16_inst_mst_rreq_ready                     : std_logic;
  signal RDAW64DW512LW8BS1BM16_inst_mst_rreq_addr                      : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_mst_rreq_len                       : std_logic_vector(BUS_LEN_WIDTH - 1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_mst_rdat_valid                     : std_logic;
  signal RDAW64DW512LW8BS1BM16_inst_mst_rdat_ready                     : std_logic;
  signal RDAW64DW512LW8BS1BM16_inst_mst_rdat_data                      : std_logic_vector(BUS_DATA_WIDTH - 1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_mst_rdat_last                      : std_logic;

  signal RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid                     : std_logic_vector(6 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready                     : std_logic_vector(6 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr                      : std_logic_vector(7 * BUS_ADDR_WIDTH - 1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len                       : std_logic_vector(7 * BUS_LEN_WIDTH - 1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid                     : std_logic_vector(6 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready                     : std_logic_vector(6 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data                      : std_logic_vector(7 * BUS_DATA_WIDTH - 1 downto 0);
  signal RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last                      : std_logic_vector(6 downto 0);

  signal WRAW64DW512LW8BS1BM16_inst_mst_wreq_valid                     : std_logic;
  signal WRAW64DW512LW8BS1BM16_inst_mst_wreq_ready                     : std_logic;
  signal WRAW64DW512LW8BS1BM16_inst_mst_wreq_addr                      : std_logic_vector(BUS_ADDR_WIDTH - 1 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_mst_wreq_len                       : std_logic_vector(BUS_LEN_WIDTH - 1 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_mst_wdat_valid                     : std_logic;
  signal WRAW64DW512LW8BS1BM16_inst_mst_wdat_ready                     : std_logic;
  signal WRAW64DW512LW8BS1BM16_inst_mst_wdat_data                      : std_logic_vector(BUS_DATA_WIDTH - 1 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_mst_wdat_strobe                    : std_logic_vector(BUS_DATA_WIDTH/8 - 1 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_mst_wdat_last                      : std_logic;

  signal WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid                     : std_logic_vector(9 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready                     : std_logic_vector(9 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr                      : std_logic_vector(10 * BUS_ADDR_WIDTH - 1 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len                       : std_logic_vector(10 * BUS_LEN_WIDTH - 1 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid                     : std_logic_vector(9 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready                     : std_logic_vector(9 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data                      : std_logic_vector(10 * BUS_DATA_WIDTH - 1 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe                    : std_logic_vector(10 * BUS_DATA_WIDTH/8 - 1 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last                      : std_logic_vector(9 downto 0);
begin
  PriceSummary_Nucleus_inst : PriceSummary_Nucleus
  generic map(
    INDEX_WIDTH                     => INDEX_WIDTH,
    TAG_WIDTH                       => TAG_WIDTH,
    L_QUANTITY_BUS_ADDR_WIDTH       => BUS_ADDR_WIDTH,
    L_EXTENDEDPRICE_BUS_ADDR_WIDTH  => BUS_ADDR_WIDTH,
    L_DISCOUNT_BUS_ADDR_WIDTH       => BUS_ADDR_WIDTH,
    L_TAX_BUS_ADDR_WIDTH            => BUS_ADDR_WIDTH,
    L_RETURNFLAG_BUS_ADDR_WIDTH     => BUS_ADDR_WIDTH,
    L_LINESTATUS_BUS_ADDR_WIDTH     => BUS_ADDR_WIDTH,
    L_SHIPDATE_BUS_ADDR_WIDTH       => BUS_ADDR_WIDTH,
    L_RETURNFLAG_O_BUS_ADDR_WIDTH   => BUS_ADDR_WIDTH,
    L_LINESTATUS_O_BUS_ADDR_WIDTH   => BUS_ADDR_WIDTH,
    L_SUM_QTY_BUS_ADDR_WIDTH        => BUS_ADDR_WIDTH,
    L_SUM_BASE_PRICE_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_SUM_DISC_PRICE_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_SUM_CHARGE_BUS_ADDR_WIDTH     => BUS_ADDR_WIDTH,
    L_AVG_QTY_BUS_ADDR_WIDTH        => BUS_ADDR_WIDTH,
    L_AVG_PRICE_BUS_ADDR_WIDTH      => BUS_ADDR_WIDTH,
    L_AVG_DISC_BUS_ADDR_WIDTH       => BUS_ADDR_WIDTH,
    L_COUNT_ORDER_BUS_ADDR_WIDTH    => BUS_ADDR_WIDTH
  )
  port map(
    kcd_clk                       => kcd_clk,
    kcd_reset                     => kcd_reset,
    mmio_awvalid                  => PriceSummary_Nucleus_inst_mmio_awvalid,
    mmio_awready                  => PriceSummary_Nucleus_inst_mmio_awready,
    mmio_awaddr                   => PriceSummary_Nucleus_inst_mmio_awaddr,
    mmio_wvalid                   => PriceSummary_Nucleus_inst_mmio_wvalid,
    mmio_wready                   => PriceSummary_Nucleus_inst_mmio_wready,
    mmio_wdata                    => PriceSummary_Nucleus_inst_mmio_wdata,
    mmio_wstrb                    => PriceSummary_Nucleus_inst_mmio_wstrb,
    mmio_bvalid                   => PriceSummary_Nucleus_inst_mmio_bvalid,
    mmio_bready                   => PriceSummary_Nucleus_inst_mmio_bready,
    mmio_bresp                    => PriceSummary_Nucleus_inst_mmio_bresp,
    mmio_arvalid                  => PriceSummary_Nucleus_inst_mmio_arvalid,
    mmio_arready                  => PriceSummary_Nucleus_inst_mmio_arready,
    mmio_araddr                   => PriceSummary_Nucleus_inst_mmio_araddr,
    mmio_rvalid                   => PriceSummary_Nucleus_inst_mmio_rvalid,
    mmio_rready                   => PriceSummary_Nucleus_inst_mmio_rready,
    mmio_rdata                    => PriceSummary_Nucleus_inst_mmio_rdata,
    mmio_rresp                    => PriceSummary_Nucleus_inst_mmio_rresp,
    l_quantity_valid              => PriceSummary_Nucleus_inst_l_quantity_valid,
    l_quantity_ready              => PriceSummary_Nucleus_inst_l_quantity_ready,
    l_quantity_dvalid             => PriceSummary_Nucleus_inst_l_quantity_dvalid,
    l_quantity_last               => PriceSummary_Nucleus_inst_l_quantity_last,
    l_quantity                    => PriceSummary_Nucleus_inst_l_quantity,
    l_extendedprice_valid         => PriceSummary_Nucleus_inst_l_extendedprice_valid,
    l_extendedprice_ready         => PriceSummary_Nucleus_inst_l_extendedprice_ready,
    l_extendedprice_dvalid        => PriceSummary_Nucleus_inst_l_extendedprice_dvalid,
    l_extendedprice_last          => PriceSummary_Nucleus_inst_l_extendedprice_last,
    l_extendedprice               => PriceSummary_Nucleus_inst_l_extendedprice,
    l_discount_valid              => PriceSummary_Nucleus_inst_l_discount_valid,
    l_discount_ready              => PriceSummary_Nucleus_inst_l_discount_ready,
    l_discount_dvalid             => PriceSummary_Nucleus_inst_l_discount_dvalid,
    l_discount_last               => PriceSummary_Nucleus_inst_l_discount_last,
    l_discount                    => PriceSummary_Nucleus_inst_l_discount,
    l_tax_valid                   => PriceSummary_Nucleus_inst_l_tax_valid,
    l_tax_ready                   => PriceSummary_Nucleus_inst_l_tax_ready,
    l_tax_dvalid                  => PriceSummary_Nucleus_inst_l_tax_dvalid,
    l_tax_last                    => PriceSummary_Nucleus_inst_l_tax_last,
    l_tax                         => PriceSummary_Nucleus_inst_l_tax,
    l_returnflag_valid            => PriceSummary_Nucleus_inst_l_returnflag_valid,
    l_returnflag_ready            => PriceSummary_Nucleus_inst_l_returnflag_ready,
    l_returnflag_dvalid           => PriceSummary_Nucleus_inst_l_returnflag_dvalid,
    l_returnflag_last             => PriceSummary_Nucleus_inst_l_returnflag_last,
    l_returnflag_length           => PriceSummary_Nucleus_inst_l_returnflag_length,
    l_returnflag_count            => PriceSummary_Nucleus_inst_l_returnflag_count,
    l_returnflag_chars_valid      => PriceSummary_Nucleus_inst_l_returnflag_chars_valid,
    l_returnflag_chars_ready      => PriceSummary_Nucleus_inst_l_returnflag_chars_ready,
    l_returnflag_chars_dvalid     => PriceSummary_Nucleus_inst_l_returnflag_chars_dvalid,
    l_returnflag_chars_last       => PriceSummary_Nucleus_inst_l_returnflag_chars_last,
    l_returnflag_chars            => PriceSummary_Nucleus_inst_l_returnflag_chars,
    l_returnflag_chars_count      => PriceSummary_Nucleus_inst_l_returnflag_chars_count,
    l_linestatus_valid            => PriceSummary_Nucleus_inst_l_linestatus_valid,
    l_linestatus_ready            => PriceSummary_Nucleus_inst_l_linestatus_ready,
    l_linestatus_dvalid           => PriceSummary_Nucleus_inst_l_linestatus_dvalid,
    l_linestatus_last             => PriceSummary_Nucleus_inst_l_linestatus_last,
    l_linestatus_length           => PriceSummary_Nucleus_inst_l_linestatus_length,
    l_linestatus_count            => PriceSummary_Nucleus_inst_l_linestatus_count,
    l_linestatus_chars_valid      => PriceSummary_Nucleus_inst_l_linestatus_chars_valid,
    l_linestatus_chars_ready      => PriceSummary_Nucleus_inst_l_linestatus_chars_ready,
    l_linestatus_chars_dvalid     => PriceSummary_Nucleus_inst_l_linestatus_chars_dvalid,
    l_linestatus_chars_last       => PriceSummary_Nucleus_inst_l_linestatus_chars_last,
    l_linestatus_chars            => PriceSummary_Nucleus_inst_l_linestatus_chars,
    l_linestatus_chars_count      => PriceSummary_Nucleus_inst_l_linestatus_chars_count,
    l_shipdate_valid              => PriceSummary_Nucleus_inst_l_shipdate_valid,
    l_shipdate_ready              => PriceSummary_Nucleus_inst_l_shipdate_ready,
    l_shipdate_dvalid             => PriceSummary_Nucleus_inst_l_shipdate_dvalid,
    l_shipdate_last               => PriceSummary_Nucleus_inst_l_shipdate_last,
    l_shipdate                    => PriceSummary_Nucleus_inst_l_shipdate,
    l_quantity_unl_valid          => PriceSummary_Nucleus_inst_l_quantity_unl_valid,
    l_quantity_unl_ready          => PriceSummary_Nucleus_inst_l_quantity_unl_ready,
    l_quantity_unl_tag            => PriceSummary_Nucleus_inst_l_quantity_unl_tag,
    l_extendedprice_unl_valid     => PriceSummary_Nucleus_inst_l_extendedprice_unl_valid,
    l_extendedprice_unl_ready     => PriceSummary_Nucleus_inst_l_extendedprice_unl_ready,
    l_extendedprice_unl_tag       => PriceSummary_Nucleus_inst_l_extendedprice_unl_tag,
    l_discount_unl_valid          => PriceSummary_Nucleus_inst_l_discount_unl_valid,
    l_discount_unl_ready          => PriceSummary_Nucleus_inst_l_discount_unl_ready,
    l_discount_unl_tag            => PriceSummary_Nucleus_inst_l_discount_unl_tag,
    l_tax_unl_valid               => PriceSummary_Nucleus_inst_l_tax_unl_valid,
    l_tax_unl_ready               => PriceSummary_Nucleus_inst_l_tax_unl_ready,
    l_tax_unl_tag                 => PriceSummary_Nucleus_inst_l_tax_unl_tag,
    l_returnflag_unl_valid        => PriceSummary_Nucleus_inst_l_returnflag_unl_valid,
    l_returnflag_unl_ready        => PriceSummary_Nucleus_inst_l_returnflag_unl_ready,
    l_returnflag_unl_tag          => PriceSummary_Nucleus_inst_l_returnflag_unl_tag,
    l_linestatus_unl_valid        => PriceSummary_Nucleus_inst_l_linestatus_unl_valid,
    l_linestatus_unl_ready        => PriceSummary_Nucleus_inst_l_linestatus_unl_ready,
    l_linestatus_unl_tag          => PriceSummary_Nucleus_inst_l_linestatus_unl_tag,
    l_shipdate_unl_valid          => PriceSummary_Nucleus_inst_l_shipdate_unl_valid,
    l_shipdate_unl_ready          => PriceSummary_Nucleus_inst_l_shipdate_unl_ready,
    l_shipdate_unl_tag            => PriceSummary_Nucleus_inst_l_shipdate_unl_tag,
    l_quantity_cmd_valid          => PriceSummary_Nucleus_inst_l_quantity_cmd_valid,
    l_quantity_cmd_ready          => PriceSummary_Nucleus_inst_l_quantity_cmd_ready,
    l_quantity_cmd_firstIdx       => PriceSummary_Nucleus_inst_l_quantity_cmd_firstIdx,
    l_quantity_cmd_lastIdx        => PriceSummary_Nucleus_inst_l_quantity_cmd_lastIdx,
    l_quantity_cmd_ctrl           => PriceSummary_Nucleus_inst_l_quantity_cmd_ctrl,
    l_quantity_cmd_tag            => PriceSummary_Nucleus_inst_l_quantity_cmd_tag,
    l_extendedprice_cmd_valid     => PriceSummary_Nucleus_inst_l_extendedprice_cmd_valid,
    l_extendedprice_cmd_ready     => PriceSummary_Nucleus_inst_l_extendedprice_cmd_ready,
    l_extendedprice_cmd_firstIdx  => PriceSummary_Nucleus_inst_l_extendedprice_cmd_firstIdx,
    l_extendedprice_cmd_lastIdx   => PriceSummary_Nucleus_inst_l_extendedprice_cmd_lastIdx,
    l_extendedprice_cmd_ctrl      => PriceSummary_Nucleus_inst_l_extendedprice_cmd_ctrl,
    l_extendedprice_cmd_tag       => PriceSummary_Nucleus_inst_l_extendedprice_cmd_tag,
    l_discount_cmd_valid          => PriceSummary_Nucleus_inst_l_discount_cmd_valid,
    l_discount_cmd_ready          => PriceSummary_Nucleus_inst_l_discount_cmd_ready,
    l_discount_cmd_firstIdx       => PriceSummary_Nucleus_inst_l_discount_cmd_firstIdx,
    l_discount_cmd_lastIdx        => PriceSummary_Nucleus_inst_l_discount_cmd_lastIdx,
    l_discount_cmd_ctrl           => PriceSummary_Nucleus_inst_l_discount_cmd_ctrl,
    l_discount_cmd_tag            => PriceSummary_Nucleus_inst_l_discount_cmd_tag,
    l_tax_cmd_valid               => PriceSummary_Nucleus_inst_l_tax_cmd_valid,
    l_tax_cmd_ready               => PriceSummary_Nucleus_inst_l_tax_cmd_ready,
    l_tax_cmd_firstIdx            => PriceSummary_Nucleus_inst_l_tax_cmd_firstIdx,
    l_tax_cmd_lastIdx             => PriceSummary_Nucleus_inst_l_tax_cmd_lastIdx,
    l_tax_cmd_ctrl                => PriceSummary_Nucleus_inst_l_tax_cmd_ctrl,
    l_tax_cmd_tag                 => PriceSummary_Nucleus_inst_l_tax_cmd_tag,
    l_returnflag_cmd_valid        => PriceSummary_Nucleus_inst_l_returnflag_cmd_valid,
    l_returnflag_cmd_ready        => PriceSummary_Nucleus_inst_l_returnflag_cmd_ready,
    l_returnflag_cmd_firstIdx     => PriceSummary_Nucleus_inst_l_returnflag_cmd_firstIdx,
    l_returnflag_cmd_lastIdx      => PriceSummary_Nucleus_inst_l_returnflag_cmd_lastIdx,
    l_returnflag_cmd_ctrl         => PriceSummary_Nucleus_inst_l_returnflag_cmd_ctrl,
    l_returnflag_cmd_tag          => PriceSummary_Nucleus_inst_l_returnflag_cmd_tag,
    l_linestatus_cmd_valid        => PriceSummary_Nucleus_inst_l_linestatus_cmd_valid,
    l_linestatus_cmd_ready        => PriceSummary_Nucleus_inst_l_linestatus_cmd_ready,
    l_linestatus_cmd_firstIdx     => PriceSummary_Nucleus_inst_l_linestatus_cmd_firstIdx,
    l_linestatus_cmd_lastIdx      => PriceSummary_Nucleus_inst_l_linestatus_cmd_lastIdx,
    l_linestatus_cmd_ctrl         => PriceSummary_Nucleus_inst_l_linestatus_cmd_ctrl,
    l_linestatus_cmd_tag          => PriceSummary_Nucleus_inst_l_linestatus_cmd_tag,
    l_shipdate_cmd_valid          => PriceSummary_Nucleus_inst_l_shipdate_cmd_valid,
    l_shipdate_cmd_ready          => PriceSummary_Nucleus_inst_l_shipdate_cmd_ready,
    l_shipdate_cmd_firstIdx       => PriceSummary_Nucleus_inst_l_shipdate_cmd_firstIdx,
    l_shipdate_cmd_lastIdx        => PriceSummary_Nucleus_inst_l_shipdate_cmd_lastIdx,
    l_shipdate_cmd_ctrl           => PriceSummary_Nucleus_inst_l_shipdate_cmd_ctrl,
    l_shipdate_cmd_tag            => PriceSummary_Nucleus_inst_l_shipdate_cmd_tag,
    l_returnflag_o_valid          => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_valid,
    l_returnflag_o_ready          => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_ready,
    l_returnflag_o_dvalid         => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_dvalid,
    l_returnflag_o_last           => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_last,
    l_returnflag_o_length         => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_length,
    l_returnflag_o_count          => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_count,
    l_returnflag_o_chars_valid    => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_valid,
    l_returnflag_o_chars_ready    => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_ready,
    l_returnflag_o_chars_dvalid   => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_dvalid,
    l_returnflag_o_chars_last     => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_last,
    l_returnflag_o_chars          => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars,
    l_returnflag_o_chars_count    => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_count,
    l_linestatus_o_valid          => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_valid,
    l_linestatus_o_ready          => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_ready,
    l_linestatus_o_dvalid         => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_dvalid,
    l_linestatus_o_last           => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_last,
    l_linestatus_o_length         => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_length,
    l_linestatus_o_count          => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_count,
    l_linestatus_o_chars_valid    => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_valid,
    l_linestatus_o_chars_ready    => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_ready,
    l_linestatus_o_chars_dvalid   => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_dvalid,
    l_linestatus_o_chars_last     => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_last,
    l_linestatus_o_chars          => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars,
    l_linestatus_o_chars_count    => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_count,
    l_sum_qty_valid               => PriceSummaryWriter_Nucleus_inst_l_sum_qty_valid,
    l_sum_qty_ready               => PriceSummaryWriter_Nucleus_inst_l_sum_qty_ready,
    l_sum_qty_dvalid              => PriceSummaryWriter_Nucleus_inst_l_sum_qty_dvalid,
    l_sum_qty_last                => PriceSummaryWriter_Nucleus_inst_l_sum_qty_last,
    l_sum_qty                     => PriceSummaryWriter_Nucleus_inst_l_sum_qty,
    l_sum_base_price_valid        => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_valid,
    l_sum_base_price_ready        => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_ready,
    l_sum_base_price_dvalid       => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_dvalid,
    l_sum_base_price_last         => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_last,
    l_sum_base_price              => PriceSummaryWriter_Nucleus_inst_l_sum_base_price,
    l_sum_disc_price_valid        => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_valid,
    l_sum_disc_price_ready        => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_ready,
    l_sum_disc_price_dvalid       => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_dvalid,
    l_sum_disc_price_last         => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_last,
    l_sum_disc_price              => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price,
    l_sum_charge_valid            => PriceSummaryWriter_Nucleus_inst_l_sum_charge_valid,
    l_sum_charge_ready            => PriceSummaryWriter_Nucleus_inst_l_sum_charge_ready,
    l_sum_charge_dvalid           => PriceSummaryWriter_Nucleus_inst_l_sum_charge_dvalid,
    l_sum_charge_last             => PriceSummaryWriter_Nucleus_inst_l_sum_charge_last,
    l_sum_charge                  => PriceSummaryWriter_Nucleus_inst_l_sum_charge,
    l_avg_qty_valid               => PriceSummaryWriter_Nucleus_inst_l_avg_qty_valid,
    l_avg_qty_ready               => PriceSummaryWriter_Nucleus_inst_l_avg_qty_ready,
    l_avg_qty_dvalid              => PriceSummaryWriter_Nucleus_inst_l_avg_qty_dvalid,
    l_avg_qty_last                => PriceSummaryWriter_Nucleus_inst_l_avg_qty_last,
    l_avg_qty                     => PriceSummaryWriter_Nucleus_inst_l_avg_qty,
    l_avg_price_valid             => PriceSummaryWriter_Nucleus_inst_l_avg_price_valid,
    l_avg_price_ready             => PriceSummaryWriter_Nucleus_inst_l_avg_price_ready,
    l_avg_price_dvalid            => PriceSummaryWriter_Nucleus_inst_l_avg_price_dvalid,
    l_avg_price_last              => PriceSummaryWriter_Nucleus_inst_l_avg_price_last,
    l_avg_price                   => PriceSummaryWriter_Nucleus_inst_l_avg_price,
    l_avg_disc_valid              => PriceSummaryWriter_Nucleus_inst_l_avg_disc_valid,
    l_avg_disc_ready              => PriceSummaryWriter_Nucleus_inst_l_avg_disc_ready,
    l_avg_disc_dvalid             => PriceSummaryWriter_Nucleus_inst_l_avg_disc_dvalid,
    l_avg_disc_last               => PriceSummaryWriter_Nucleus_inst_l_avg_disc_last,
    l_avg_disc                    => PriceSummaryWriter_Nucleus_inst_l_avg_disc,
    l_count_order_valid           => PriceSummaryWriter_Nucleus_inst_l_count_order_valid,
    l_count_order_ready           => PriceSummaryWriter_Nucleus_inst_l_count_order_ready,
    l_count_order_dvalid          => PriceSummaryWriter_Nucleus_inst_l_count_order_dvalid,
    l_count_order_last            => PriceSummaryWriter_Nucleus_inst_l_count_order_last,
    l_count_order                 => PriceSummaryWriter_Nucleus_inst_l_count_order,
    l_returnflag_o_unl_valid      => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_unl_valid,
    l_returnflag_o_unl_ready      => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_unl_ready,
    l_returnflag_o_unl_tag        => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_unl_tag,
    l_linestatus_o_unl_valid      => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_unl_valid,
    l_linestatus_o_unl_ready      => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_unl_ready,
    l_linestatus_o_unl_tag        => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_unl_tag,
    l_sum_qty_unl_valid           => PriceSummaryWriter_Nucleus_inst_l_sum_qty_unl_valid,
    l_sum_qty_unl_ready           => PriceSummaryWriter_Nucleus_inst_l_sum_qty_unl_ready,
    l_sum_qty_unl_tag             => PriceSummaryWriter_Nucleus_inst_l_sum_qty_unl_tag,
    l_sum_base_price_unl_valid    => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_unl_valid,
    l_sum_base_price_unl_ready    => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_unl_ready,
    l_sum_base_price_unl_tag      => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_unl_tag,
    l_sum_disc_price_unl_valid    => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_unl_valid,
    l_sum_disc_price_unl_ready    => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_unl_ready,
    l_sum_disc_price_unl_tag      => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_unl_tag,
    l_sum_charge_unl_valid        => PriceSummaryWriter_Nucleus_inst_l_sum_charge_unl_valid,
    l_sum_charge_unl_ready        => PriceSummaryWriter_Nucleus_inst_l_sum_charge_unl_ready,
    l_sum_charge_unl_tag          => PriceSummaryWriter_Nucleus_inst_l_sum_charge_unl_tag,
    l_avg_qty_unl_valid           => PriceSummaryWriter_Nucleus_inst_l_avg_qty_unl_valid,
    l_avg_qty_unl_ready           => PriceSummaryWriter_Nucleus_inst_l_avg_qty_unl_ready,
    l_avg_qty_unl_tag             => PriceSummaryWriter_Nucleus_inst_l_avg_qty_unl_tag,
    l_avg_price_unl_valid         => PriceSummaryWriter_Nucleus_inst_l_avg_price_unl_valid,
    l_avg_price_unl_ready         => PriceSummaryWriter_Nucleus_inst_l_avg_price_unl_ready,
    l_avg_price_unl_tag           => PriceSummaryWriter_Nucleus_inst_l_avg_price_unl_tag,
    l_avg_disc_unl_valid          => PriceSummaryWriter_Nucleus_inst_l_avg_disc_unl_valid,
    l_avg_disc_unl_ready          => PriceSummaryWriter_Nucleus_inst_l_avg_disc_unl_ready,
    l_avg_disc_unl_tag            => PriceSummaryWriter_Nucleus_inst_l_avg_disc_unl_tag,
    l_count_order_unl_valid       => PriceSummaryWriter_Nucleus_inst_l_count_order_unl_valid,
    l_count_order_unl_ready       => PriceSummaryWriter_Nucleus_inst_l_count_order_unl_ready,
    l_count_order_unl_tag         => PriceSummaryWriter_Nucleus_inst_l_count_order_unl_tag,
    l_returnflag_o_cmd_valid      => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_valid,
    l_returnflag_o_cmd_ready      => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_ready,
    l_returnflag_o_cmd_firstIdx   => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_firstIdx,
    l_returnflag_o_cmd_lastIdx    => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_lastIdx,
    l_returnflag_o_cmd_ctrl       => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_ctrl,
    l_returnflag_o_cmd_tag        => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_tag,
    l_linestatus_o_cmd_valid      => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_valid,
    l_linestatus_o_cmd_ready      => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_ready,
    l_linestatus_o_cmd_firstIdx   => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_firstIdx,
    l_linestatus_o_cmd_lastIdx    => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_lastIdx,
    l_linestatus_o_cmd_ctrl       => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_ctrl,
    l_linestatus_o_cmd_tag        => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_tag,
    l_sum_qty_cmd_valid           => PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_valid,
    l_sum_qty_cmd_ready           => PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_ready,
    l_sum_qty_cmd_firstIdx        => PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_firstIdx,
    l_sum_qty_cmd_lastIdx         => PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_lastIdx,
    l_sum_qty_cmd_ctrl            => PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_ctrl,
    l_sum_qty_cmd_tag             => PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_tag,
    l_sum_base_price_cmd_valid    => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_valid,
    l_sum_base_price_cmd_ready    => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_ready,
    l_sum_base_price_cmd_firstIdx => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_firstIdx,
    l_sum_base_price_cmd_lastIdx  => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_lastIdx,
    l_sum_base_price_cmd_ctrl     => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_ctrl,
    l_sum_base_price_cmd_tag      => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_tag,
    l_sum_disc_price_cmd_valid    => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_valid,
    l_sum_disc_price_cmd_ready    => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_ready,
    l_sum_disc_price_cmd_firstIdx => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_firstIdx,
    l_sum_disc_price_cmd_lastIdx  => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_lastIdx,
    l_sum_disc_price_cmd_ctrl     => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_ctrl,
    l_sum_disc_price_cmd_tag      => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_tag,
    l_sum_charge_cmd_valid        => PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_valid,
    l_sum_charge_cmd_ready        => PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_ready,
    l_sum_charge_cmd_firstIdx     => PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_firstIdx,
    l_sum_charge_cmd_lastIdx      => PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_lastIdx,
    l_sum_charge_cmd_ctrl         => PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_ctrl,
    l_sum_charge_cmd_tag          => PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_tag,
    l_avg_qty_cmd_valid           => PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_valid,
    l_avg_qty_cmd_ready           => PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_ready,
    l_avg_qty_cmd_firstIdx        => PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_firstIdx,
    l_avg_qty_cmd_lastIdx         => PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_lastIdx,
    l_avg_qty_cmd_ctrl            => PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_ctrl,
    l_avg_qty_cmd_tag             => PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_tag,
    l_avg_price_cmd_valid         => PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_valid,
    l_avg_price_cmd_ready         => PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_ready,
    l_avg_price_cmd_firstIdx      => PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_firstIdx,
    l_avg_price_cmd_lastIdx       => PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_lastIdx,
    l_avg_price_cmd_ctrl          => PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_ctrl,
    l_avg_price_cmd_tag           => PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_tag,
    l_avg_disc_cmd_valid          => PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_valid,
    l_avg_disc_cmd_ready          => PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_ready,
    l_avg_disc_cmd_firstIdx       => PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_firstIdx,
    l_avg_disc_cmd_lastIdx        => PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_lastIdx,
    l_avg_disc_cmd_ctrl           => PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_ctrl,
    l_avg_disc_cmd_tag            => PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_tag,
    l_count_order_cmd_valid       => PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_valid,
    l_count_order_cmd_ready       => PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_ready,
    l_count_order_cmd_firstIdx    => PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_firstIdx,
    l_count_order_cmd_lastIdx     => PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_lastIdx,
    l_count_order_cmd_ctrl        => PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_ctrl,
    l_count_order_cmd_tag         => PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_tag
  );

  PriceSummary_l_inst : PriceSummary_l
  generic map(
    INDEX_WIDTH                         => INDEX_WIDTH,
    TAG_WIDTH                           => TAG_WIDTH,
    L_QUANTITY_BUS_ADDR_WIDTH           => BUS_ADDR_WIDTH,
    L_QUANTITY_BUS_DATA_WIDTH           => BUS_DATA_WIDTH,
    L_QUANTITY_BUS_LEN_WIDTH            => BUS_LEN_WIDTH,
    L_QUANTITY_BUS_BURST_STEP_LEN       => BUS_BURST_STEP_LEN,
    L_QUANTITY_BUS_BURST_MAX_LEN        => BUS_BURST_MAX_LEN,
    L_EXTENDEDPRICE_BUS_ADDR_WIDTH      => BUS_ADDR_WIDTH,
    L_EXTENDEDPRICE_BUS_DATA_WIDTH      => BUS_DATA_WIDTH,
    L_EXTENDEDPRICE_BUS_LEN_WIDTH       => BUS_LEN_WIDTH,
    L_EXTENDEDPRICE_BUS_BURST_STEP_LEN  => BUS_BURST_STEP_LEN,
    L_EXTENDEDPRICE_BUS_BURST_MAX_LEN   => BUS_BURST_MAX_LEN,
    L_DISCOUNT_BUS_ADDR_WIDTH           => BUS_ADDR_WIDTH,
    L_DISCOUNT_BUS_DATA_WIDTH           => BUS_DATA_WIDTH,
    L_DISCOUNT_BUS_LEN_WIDTH            => BUS_LEN_WIDTH,
    L_DISCOUNT_BUS_BURST_STEP_LEN       => BUS_BURST_STEP_LEN,
    L_DISCOUNT_BUS_BURST_MAX_LEN        => BUS_BURST_MAX_LEN,
    L_TAX_BUS_ADDR_WIDTH                => BUS_ADDR_WIDTH,
    L_TAX_BUS_DATA_WIDTH                => BUS_DATA_WIDTH,
    L_TAX_BUS_LEN_WIDTH                 => BUS_LEN_WIDTH,
    L_TAX_BUS_BURST_STEP_LEN            => BUS_BURST_STEP_LEN,
    L_TAX_BUS_BURST_MAX_LEN             => BUS_BURST_MAX_LEN,
    L_RETURNFLAG_BUS_ADDR_WIDTH         => BUS_ADDR_WIDTH,
    L_RETURNFLAG_BUS_DATA_WIDTH         => BUS_DATA_WIDTH,
    L_RETURNFLAG_BUS_LEN_WIDTH          => BUS_LEN_WIDTH,
    L_RETURNFLAG_BUS_BURST_STEP_LEN     => BUS_BURST_STEP_LEN,
    L_RETURNFLAG_BUS_BURST_MAX_LEN      => BUS_BURST_MAX_LEN,
    L_LINESTATUS_BUS_ADDR_WIDTH         => BUS_ADDR_WIDTH,
    L_LINESTATUS_BUS_DATA_WIDTH         => BUS_DATA_WIDTH,
    L_LINESTATUS_BUS_LEN_WIDTH          => BUS_LEN_WIDTH,
    L_LINESTATUS_BUS_BURST_STEP_LEN     => BUS_BURST_STEP_LEN,
    L_LINESTATUS_BUS_BURST_MAX_LEN      => BUS_BURST_MAX_LEN,
    L_SHIPDATE_BUS_ADDR_WIDTH           => BUS_ADDR_WIDTH,
    L_SHIPDATE_BUS_DATA_WIDTH           => BUS_DATA_WIDTH,
    L_SHIPDATE_BUS_LEN_WIDTH            => BUS_LEN_WIDTH,
    L_SHIPDATE_BUS_BURST_STEP_LEN       => BUS_BURST_STEP_LEN,
    L_SHIPDATE_BUS_BURST_MAX_LEN        => BUS_BURST_MAX_LEN,
    L_RETURNFLAG_O_BUS_ADDR_WIDTH       => BUS_ADDR_WIDTH,
    L_RETURNFLAG_O_BUS_DATA_WIDTH       => BUS_DATA_WIDTH,
    L_RETURNFLAG_O_BUS_LEN_WIDTH        => BUS_LEN_WIDTH,
    L_RETURNFLAG_O_BUS_BURST_STEP_LEN   => BUS_BURST_STEP_LEN,
    L_RETURNFLAG_O_BUS_BURST_MAX_LEN    => BUS_BURST_MAX_LEN,
    L_LINESTATUS_O_BUS_ADDR_WIDTH       => BUS_ADDR_WIDTH,
    L_LINESTATUS_O_BUS_DATA_WIDTH       => BUS_DATA_WIDTH,
    L_LINESTATUS_O_BUS_LEN_WIDTH        => BUS_LEN_WIDTH,
    L_LINESTATUS_O_BUS_BURST_STEP_LEN   => BUS_BURST_STEP_LEN,
    L_LINESTATUS_O_BUS_BURST_MAX_LEN    => BUS_BURST_MAX_LEN,
    L_SUM_QTY_BUS_ADDR_WIDTH            => BUS_ADDR_WIDTH,
    L_SUM_QTY_BUS_DATA_WIDTH            => BUS_DATA_WIDTH,
    L_SUM_QTY_BUS_LEN_WIDTH             => BUS_LEN_WIDTH,
    L_SUM_QTY_BUS_BURST_STEP_LEN        => BUS_BURST_STEP_LEN,
    L_SUM_QTY_BUS_BURST_MAX_LEN         => BUS_BURST_MAX_LEN,
    L_SUM_BASE_PRICE_BUS_ADDR_WIDTH     => BUS_ADDR_WIDTH,
    L_SUM_BASE_PRICE_BUS_DATA_WIDTH     => BUS_DATA_WIDTH,
    L_SUM_BASE_PRICE_BUS_LEN_WIDTH      => BUS_LEN_WIDTH,
    L_SUM_BASE_PRICE_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
    L_SUM_BASE_PRICE_BUS_BURST_MAX_LEN  => BUS_BURST_MAX_LEN,
    L_SUM_DISC_PRICE_BUS_ADDR_WIDTH     => BUS_ADDR_WIDTH,
    L_SUM_DISC_PRICE_BUS_DATA_WIDTH     => BUS_DATA_WIDTH,
    L_SUM_DISC_PRICE_BUS_LEN_WIDTH      => BUS_LEN_WIDTH,
    L_SUM_DISC_PRICE_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
    L_SUM_DISC_PRICE_BUS_BURST_MAX_LEN  => BUS_BURST_MAX_LEN,
    L_SUM_CHARGE_BUS_ADDR_WIDTH         => BUS_ADDR_WIDTH,
    L_SUM_CHARGE_BUS_DATA_WIDTH         => BUS_DATA_WIDTH,
    L_SUM_CHARGE_BUS_LEN_WIDTH          => BUS_LEN_WIDTH,
    L_SUM_CHARGE_BUS_BURST_STEP_LEN     => BUS_BURST_STEP_LEN,
    L_SUM_CHARGE_BUS_BURST_MAX_LEN      => BUS_BURST_MAX_LEN,
    L_AVG_QTY_BUS_ADDR_WIDTH            => BUS_ADDR_WIDTH,
    L_AVG_QTY_BUS_DATA_WIDTH            => BUS_DATA_WIDTH,
    L_AVG_QTY_BUS_LEN_WIDTH             => BUS_LEN_WIDTH,
    L_AVG_QTY_BUS_BURST_STEP_LEN        => BUS_BURST_STEP_LEN,
    L_AVG_QTY_BUS_BURST_MAX_LEN         => BUS_BURST_MAX_LEN,
    L_AVG_PRICE_BUS_ADDR_WIDTH          => BUS_ADDR_WIDTH,
    L_AVG_PRICE_BUS_DATA_WIDTH          => BUS_DATA_WIDTH,
    L_AVG_PRICE_BUS_LEN_WIDTH           => BUS_LEN_WIDTH,
    L_AVG_PRICE_BUS_BURST_STEP_LEN      => BUS_BURST_STEP_LEN,
    L_AVG_PRICE_BUS_BURST_MAX_LEN       => BUS_BURST_MAX_LEN,
    L_AVG_DISC_BUS_ADDR_WIDTH           => BUS_ADDR_WIDTH,
    L_AVG_DISC_BUS_DATA_WIDTH           => BUS_DATA_WIDTH,
    L_AVG_DISC_BUS_LEN_WIDTH            => BUS_LEN_WIDTH,
    L_AVG_DISC_BUS_BURST_STEP_LEN       => BUS_BURST_STEP_LEN,
    L_AVG_DISC_BUS_BURST_MAX_LEN        => BUS_BURST_MAX_LEN,
    L_COUNT_ORDER_BUS_ADDR_WIDTH        => BUS_ADDR_WIDTH,
    L_COUNT_ORDER_BUS_DATA_WIDTH        => BUS_DATA_WIDTH,
    L_COUNT_ORDER_BUS_LEN_WIDTH         => BUS_LEN_WIDTH,
    L_COUNT_ORDER_BUS_BURST_STEP_LEN    => BUS_BURST_STEP_LEN,
    L_COUNT_ORDER_BUS_BURST_MAX_LEN     => BUS_BURST_MAX_LEN
  )
  port map(
    bcd_clk                          => bcd_clk,
    bcd_reset                        => bcd_reset,
    kcd_clk                          => kcd_clk,
    kcd_reset                        => kcd_reset,
    l_quantity_valid                 => PriceSummary_l_inst_l_quantity_valid,
    l_quantity_ready                 => PriceSummary_l_inst_l_quantity_ready,
    l_quantity_dvalid                => PriceSummary_l_inst_l_quantity_dvalid,
    l_quantity_last                  => PriceSummary_l_inst_l_quantity_last,
    l_quantity                       => PriceSummary_l_inst_l_quantity,
    l_quantity_bus_rreq_valid        => PriceSummary_l_inst_l_quantity_bus_rreq_valid,
    l_quantity_bus_rreq_ready        => PriceSummary_l_inst_l_quantity_bus_rreq_ready,
    l_quantity_bus_rreq_addr         => PriceSummary_l_inst_l_quantity_bus_rreq_addr,
    l_quantity_bus_rreq_len          => PriceSummary_l_inst_l_quantity_bus_rreq_len,
    l_quantity_bus_rdat_valid        => PriceSummary_l_inst_l_quantity_bus_rdat_valid,
    l_quantity_bus_rdat_ready        => PriceSummary_l_inst_l_quantity_bus_rdat_ready,
    l_quantity_bus_rdat_data         => PriceSummary_l_inst_l_quantity_bus_rdat_data,
    l_quantity_bus_rdat_last         => PriceSummary_l_inst_l_quantity_bus_rdat_last,
    l_quantity_cmd_valid             => PriceSummary_l_inst_l_quantity_cmd_valid,
    l_quantity_cmd_ready             => PriceSummary_l_inst_l_quantity_cmd_ready,
    l_quantity_cmd_firstIdx          => PriceSummary_l_inst_l_quantity_cmd_firstIdx,
    l_quantity_cmd_lastIdx           => PriceSummary_l_inst_l_quantity_cmd_lastIdx,
    l_quantity_cmd_ctrl              => PriceSummary_l_inst_l_quantity_cmd_ctrl,
    l_quantity_cmd_tag               => PriceSummary_l_inst_l_quantity_cmd_tag,
    l_quantity_unl_valid             => PriceSummary_l_inst_l_quantity_unl_valid,
    l_quantity_unl_ready             => PriceSummary_l_inst_l_quantity_unl_ready,
    l_quantity_unl_tag               => PriceSummary_l_inst_l_quantity_unl_tag,
    l_extendedprice_valid            => PriceSummary_l_inst_l_extendedprice_valid,
    l_extendedprice_ready            => PriceSummary_l_inst_l_extendedprice_ready,
    l_extendedprice_dvalid           => PriceSummary_l_inst_l_extendedprice_dvalid,
    l_extendedprice_last             => PriceSummary_l_inst_l_extendedprice_last,
    l_extendedprice                  => PriceSummary_l_inst_l_extendedprice,
    l_extendedprice_bus_rreq_valid   => PriceSummary_l_inst_l_extendedprice_bus_rreq_valid,
    l_extendedprice_bus_rreq_ready   => PriceSummary_l_inst_l_extendedprice_bus_rreq_ready,
    l_extendedprice_bus_rreq_addr    => PriceSummary_l_inst_l_extendedprice_bus_rreq_addr,
    l_extendedprice_bus_rreq_len     => PriceSummary_l_inst_l_extendedprice_bus_rreq_len,
    l_extendedprice_bus_rdat_valid   => PriceSummary_l_inst_l_extendedprice_bus_rdat_valid,
    l_extendedprice_bus_rdat_ready   => PriceSummary_l_inst_l_extendedprice_bus_rdat_ready,
    l_extendedprice_bus_rdat_data    => PriceSummary_l_inst_l_extendedprice_bus_rdat_data,
    l_extendedprice_bus_rdat_last    => PriceSummary_l_inst_l_extendedprice_bus_rdat_last,
    l_extendedprice_cmd_valid        => PriceSummary_l_inst_l_extendedprice_cmd_valid,
    l_extendedprice_cmd_ready        => PriceSummary_l_inst_l_extendedprice_cmd_ready,
    l_extendedprice_cmd_firstIdx     => PriceSummary_l_inst_l_extendedprice_cmd_firstIdx,
    l_extendedprice_cmd_lastIdx      => PriceSummary_l_inst_l_extendedprice_cmd_lastIdx,
    l_extendedprice_cmd_ctrl         => PriceSummary_l_inst_l_extendedprice_cmd_ctrl,
    l_extendedprice_cmd_tag          => PriceSummary_l_inst_l_extendedprice_cmd_tag,
    l_extendedprice_unl_valid        => PriceSummary_l_inst_l_extendedprice_unl_valid,
    l_extendedprice_unl_ready        => PriceSummary_l_inst_l_extendedprice_unl_ready,
    l_extendedprice_unl_tag          => PriceSummary_l_inst_l_extendedprice_unl_tag,
    l_discount_valid                 => PriceSummary_l_inst_l_discount_valid,
    l_discount_ready                 => PriceSummary_l_inst_l_discount_ready,
    l_discount_dvalid                => PriceSummary_l_inst_l_discount_dvalid,
    l_discount_last                  => PriceSummary_l_inst_l_discount_last,
    l_discount                       => PriceSummary_l_inst_l_discount,
    l_discount_bus_rreq_valid        => PriceSummary_l_inst_l_discount_bus_rreq_valid,
    l_discount_bus_rreq_ready        => PriceSummary_l_inst_l_discount_bus_rreq_ready,
    l_discount_bus_rreq_addr         => PriceSummary_l_inst_l_discount_bus_rreq_addr,
    l_discount_bus_rreq_len          => PriceSummary_l_inst_l_discount_bus_rreq_len,
    l_discount_bus_rdat_valid        => PriceSummary_l_inst_l_discount_bus_rdat_valid,
    l_discount_bus_rdat_ready        => PriceSummary_l_inst_l_discount_bus_rdat_ready,
    l_discount_bus_rdat_data         => PriceSummary_l_inst_l_discount_bus_rdat_data,
    l_discount_bus_rdat_last         => PriceSummary_l_inst_l_discount_bus_rdat_last,
    l_discount_cmd_valid             => PriceSummary_l_inst_l_discount_cmd_valid,
    l_discount_cmd_ready             => PriceSummary_l_inst_l_discount_cmd_ready,
    l_discount_cmd_firstIdx          => PriceSummary_l_inst_l_discount_cmd_firstIdx,
    l_discount_cmd_lastIdx           => PriceSummary_l_inst_l_discount_cmd_lastIdx,
    l_discount_cmd_ctrl              => PriceSummary_l_inst_l_discount_cmd_ctrl,
    l_discount_cmd_tag               => PriceSummary_l_inst_l_discount_cmd_tag,
    l_discount_unl_valid             => PriceSummary_l_inst_l_discount_unl_valid,
    l_discount_unl_ready             => PriceSummary_l_inst_l_discount_unl_ready,
    l_discount_unl_tag               => PriceSummary_l_inst_l_discount_unl_tag,
    l_tax_valid                      => PriceSummary_l_inst_l_tax_valid,
    l_tax_ready                      => PriceSummary_l_inst_l_tax_ready,
    l_tax_dvalid                     => PriceSummary_l_inst_l_tax_dvalid,
    l_tax_last                       => PriceSummary_l_inst_l_tax_last,
    l_tax                            => PriceSummary_l_inst_l_tax,
    l_tax_bus_rreq_valid             => PriceSummary_l_inst_l_tax_bus_rreq_valid,
    l_tax_bus_rreq_ready             => PriceSummary_l_inst_l_tax_bus_rreq_ready,
    l_tax_bus_rreq_addr              => PriceSummary_l_inst_l_tax_bus_rreq_addr,
    l_tax_bus_rreq_len               => PriceSummary_l_inst_l_tax_bus_rreq_len,
    l_tax_bus_rdat_valid             => PriceSummary_l_inst_l_tax_bus_rdat_valid,
    l_tax_bus_rdat_ready             => PriceSummary_l_inst_l_tax_bus_rdat_ready,
    l_tax_bus_rdat_data              => PriceSummary_l_inst_l_tax_bus_rdat_data,
    l_tax_bus_rdat_last              => PriceSummary_l_inst_l_tax_bus_rdat_last,
    l_tax_cmd_valid                  => PriceSummary_l_inst_l_tax_cmd_valid,
    l_tax_cmd_ready                  => PriceSummary_l_inst_l_tax_cmd_ready,
    l_tax_cmd_firstIdx               => PriceSummary_l_inst_l_tax_cmd_firstIdx,
    l_tax_cmd_lastIdx                => PriceSummary_l_inst_l_tax_cmd_lastIdx,
    l_tax_cmd_ctrl                   => PriceSummary_l_inst_l_tax_cmd_ctrl,
    l_tax_cmd_tag                    => PriceSummary_l_inst_l_tax_cmd_tag,
    l_tax_unl_valid                  => PriceSummary_l_inst_l_tax_unl_valid,
    l_tax_unl_ready                  => PriceSummary_l_inst_l_tax_unl_ready,
    l_tax_unl_tag                    => PriceSummary_l_inst_l_tax_unl_tag,
    l_returnflag_valid               => PriceSummary_l_inst_l_returnflag_valid,
    l_returnflag_ready               => PriceSummary_l_inst_l_returnflag_ready,
    l_returnflag_dvalid              => PriceSummary_l_inst_l_returnflag_dvalid,
    l_returnflag_last                => PriceSummary_l_inst_l_returnflag_last,
    l_returnflag_length              => PriceSummary_l_inst_l_returnflag_length,
    l_returnflag_count               => PriceSummary_l_inst_l_returnflag_count,
    l_returnflag_chars_valid         => PriceSummary_l_inst_l_returnflag_chars_valid,
    l_returnflag_chars_ready         => PriceSummary_l_inst_l_returnflag_chars_ready,
    l_returnflag_chars_dvalid        => PriceSummary_l_inst_l_returnflag_chars_dvalid,
    l_returnflag_chars_last          => PriceSummary_l_inst_l_returnflag_chars_last,
    l_returnflag_chars               => PriceSummary_l_inst_l_returnflag_chars,
    l_returnflag_chars_count         => PriceSummary_l_inst_l_returnflag_chars_count,
    l_returnflag_bus_rreq_valid      => PriceSummary_l_inst_l_returnflag_bus_rreq_valid,
    l_returnflag_bus_rreq_ready      => PriceSummary_l_inst_l_returnflag_bus_rreq_ready,
    l_returnflag_bus_rreq_addr       => PriceSummary_l_inst_l_returnflag_bus_rreq_addr,
    l_returnflag_bus_rreq_len        => PriceSummary_l_inst_l_returnflag_bus_rreq_len,
    l_returnflag_bus_rdat_valid      => PriceSummary_l_inst_l_returnflag_bus_rdat_valid,
    l_returnflag_bus_rdat_ready      => PriceSummary_l_inst_l_returnflag_bus_rdat_ready,
    l_returnflag_bus_rdat_data       => PriceSummary_l_inst_l_returnflag_bus_rdat_data,
    l_returnflag_bus_rdat_last       => PriceSummary_l_inst_l_returnflag_bus_rdat_last,
    l_returnflag_cmd_valid           => PriceSummary_l_inst_l_returnflag_cmd_valid,
    l_returnflag_cmd_ready           => PriceSummary_l_inst_l_returnflag_cmd_ready,
    l_returnflag_cmd_firstIdx        => PriceSummary_l_inst_l_returnflag_cmd_firstIdx,
    l_returnflag_cmd_lastIdx         => PriceSummary_l_inst_l_returnflag_cmd_lastIdx,
    l_returnflag_cmd_ctrl            => PriceSummary_l_inst_l_returnflag_cmd_ctrl,
    l_returnflag_cmd_tag             => PriceSummary_l_inst_l_returnflag_cmd_tag,
    l_returnflag_unl_valid           => PriceSummary_l_inst_l_returnflag_unl_valid,
    l_returnflag_unl_ready           => PriceSummary_l_inst_l_returnflag_unl_ready,
    l_returnflag_unl_tag             => PriceSummary_l_inst_l_returnflag_unl_tag,
    l_linestatus_valid               => PriceSummary_l_inst_l_linestatus_valid,
    l_linestatus_ready               => PriceSummary_l_inst_l_linestatus_ready,
    l_linestatus_dvalid              => PriceSummary_l_inst_l_linestatus_dvalid,
    l_linestatus_last                => PriceSummary_l_inst_l_linestatus_last,
    l_linestatus_length              => PriceSummary_l_inst_l_linestatus_length,
    l_linestatus_count               => PriceSummary_l_inst_l_linestatus_count,
    l_linestatus_chars_valid         => PriceSummary_l_inst_l_linestatus_chars_valid,
    l_linestatus_chars_ready         => PriceSummary_l_inst_l_linestatus_chars_ready,
    l_linestatus_chars_dvalid        => PriceSummary_l_inst_l_linestatus_chars_dvalid,
    l_linestatus_chars_last          => PriceSummary_l_inst_l_linestatus_chars_last,
    l_linestatus_chars               => PriceSummary_l_inst_l_linestatus_chars,
    l_linestatus_chars_count         => PriceSummary_l_inst_l_linestatus_chars_count,
    l_linestatus_bus_rreq_valid      => PriceSummary_l_inst_l_linestatus_bus_rreq_valid,
    l_linestatus_bus_rreq_ready      => PriceSummary_l_inst_l_linestatus_bus_rreq_ready,
    l_linestatus_bus_rreq_addr       => PriceSummary_l_inst_l_linestatus_bus_rreq_addr,
    l_linestatus_bus_rreq_len        => PriceSummary_l_inst_l_linestatus_bus_rreq_len,
    l_linestatus_bus_rdat_valid      => PriceSummary_l_inst_l_linestatus_bus_rdat_valid,
    l_linestatus_bus_rdat_ready      => PriceSummary_l_inst_l_linestatus_bus_rdat_ready,
    l_linestatus_bus_rdat_data       => PriceSummary_l_inst_l_linestatus_bus_rdat_data,
    l_linestatus_bus_rdat_last       => PriceSummary_l_inst_l_linestatus_bus_rdat_last,
    l_linestatus_cmd_valid           => PriceSummary_l_inst_l_linestatus_cmd_valid,
    l_linestatus_cmd_ready           => PriceSummary_l_inst_l_linestatus_cmd_ready,
    l_linestatus_cmd_firstIdx        => PriceSummary_l_inst_l_linestatus_cmd_firstIdx,
    l_linestatus_cmd_lastIdx         => PriceSummary_l_inst_l_linestatus_cmd_lastIdx,
    l_linestatus_cmd_ctrl            => PriceSummary_l_inst_l_linestatus_cmd_ctrl,
    l_linestatus_cmd_tag             => PriceSummary_l_inst_l_linestatus_cmd_tag,
    l_linestatus_unl_valid           => PriceSummary_l_inst_l_linestatus_unl_valid,
    l_linestatus_unl_ready           => PriceSummary_l_inst_l_linestatus_unl_ready,
    l_linestatus_unl_tag             => PriceSummary_l_inst_l_linestatus_unl_tag,
    l_shipdate_valid                 => PriceSummary_l_inst_l_shipdate_valid,
    l_shipdate_ready                 => PriceSummary_l_inst_l_shipdate_ready,
    l_shipdate_dvalid                => PriceSummary_l_inst_l_shipdate_dvalid,
    l_shipdate_last                  => PriceSummary_l_inst_l_shipdate_last,
    l_shipdate                       => PriceSummary_l_inst_l_shipdate,
    l_shipdate_bus_rreq_valid        => PriceSummary_l_inst_l_shipdate_bus_rreq_valid,
    l_shipdate_bus_rreq_ready        => PriceSummary_l_inst_l_shipdate_bus_rreq_ready,
    l_shipdate_bus_rreq_addr         => PriceSummary_l_inst_l_shipdate_bus_rreq_addr,
    l_shipdate_bus_rreq_len          => PriceSummary_l_inst_l_shipdate_bus_rreq_len,
    l_shipdate_bus_rdat_valid        => PriceSummary_l_inst_l_shipdate_bus_rdat_valid,
    l_shipdate_bus_rdat_ready        => PriceSummary_l_inst_l_shipdate_bus_rdat_ready,
    l_shipdate_bus_rdat_data         => PriceSummary_l_inst_l_shipdate_bus_rdat_data,
    l_shipdate_bus_rdat_last         => PriceSummary_l_inst_l_shipdate_bus_rdat_last,
    l_shipdate_cmd_valid             => PriceSummary_l_inst_l_shipdate_cmd_valid,
    l_shipdate_cmd_ready             => PriceSummary_l_inst_l_shipdate_cmd_ready,
    l_shipdate_cmd_firstIdx          => PriceSummary_l_inst_l_shipdate_cmd_firstIdx,
    l_shipdate_cmd_lastIdx           => PriceSummary_l_inst_l_shipdate_cmd_lastIdx,
    l_shipdate_cmd_ctrl              => PriceSummary_l_inst_l_shipdate_cmd_ctrl,
    l_shipdate_cmd_tag               => PriceSummary_l_inst_l_shipdate_cmd_tag,
    l_shipdate_unl_valid             => PriceSummary_l_inst_l_shipdate_unl_valid,
    l_shipdate_unl_ready             => PriceSummary_l_inst_l_shipdate_unl_ready,
    l_shipdate_unl_tag               => PriceSummary_l_inst_l_shipdate_unl_tag,
    l_returnflag_o_valid             => PriceSummaryWriter_l_inst_l_returnflag_o_valid,
    l_returnflag_o_ready             => PriceSummaryWriter_l_inst_l_returnflag_o_ready,
    l_returnflag_o_dvalid            => PriceSummaryWriter_l_inst_l_returnflag_o_dvalid,
    l_returnflag_o_last              => PriceSummaryWriter_l_inst_l_returnflag_o_last,
    l_returnflag_o_length            => PriceSummaryWriter_l_inst_l_returnflag_o_length,
    l_returnflag_o_count             => PriceSummaryWriter_l_inst_l_returnflag_o_count,
    l_returnflag_o_chars_valid       => PriceSummaryWriter_l_inst_l_returnflag_o_chars_valid,
    l_returnflag_o_chars_ready       => PriceSummaryWriter_l_inst_l_returnflag_o_chars_ready,
    l_returnflag_o_chars_dvalid      => PriceSummaryWriter_l_inst_l_returnflag_o_chars_dvalid,
    l_returnflag_o_chars_last        => PriceSummaryWriter_l_inst_l_returnflag_o_chars_last,
    l_returnflag_o_chars             => PriceSummaryWriter_l_inst_l_returnflag_o_chars,
    l_returnflag_o_chars_count       => PriceSummaryWriter_l_inst_l_returnflag_o_chars_count,
    l_returnflag_o_bus_wreq_valid    => PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_valid,
    l_returnflag_o_bus_wreq_ready    => PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_ready,
    l_returnflag_o_bus_wreq_addr     => PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_addr,
    l_returnflag_o_bus_wreq_len      => PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_len,
    l_returnflag_o_bus_wdat_valid    => PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_valid,
    l_returnflag_o_bus_wdat_ready    => PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_ready,
    l_returnflag_o_bus_wdat_data     => PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_data,
    l_returnflag_o_bus_wdat_strobe   => PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_strobe,
    l_returnflag_o_bus_wdat_last     => PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_last,
    l_returnflag_o_cmd_valid         => PriceSummaryWriter_l_inst_l_returnflag_o_cmd_valid,
    l_returnflag_o_cmd_ready         => PriceSummaryWriter_l_inst_l_returnflag_o_cmd_ready,
    l_returnflag_o_cmd_firstIdx      => PriceSummaryWriter_l_inst_l_returnflag_o_cmd_firstIdx,
    l_returnflag_o_cmd_lastIdx       => PriceSummaryWriter_l_inst_l_returnflag_o_cmd_lastIdx,
    l_returnflag_o_cmd_ctrl          => PriceSummaryWriter_l_inst_l_returnflag_o_cmd_ctrl,
    l_returnflag_o_cmd_tag           => PriceSummaryWriter_l_inst_l_returnflag_o_cmd_tag,
    l_returnflag_o_unl_valid         => PriceSummaryWriter_l_inst_l_returnflag_o_unl_valid,
    l_returnflag_o_unl_ready         => PriceSummaryWriter_l_inst_l_returnflag_o_unl_ready,
    l_returnflag_o_unl_tag           => PriceSummaryWriter_l_inst_l_returnflag_o_unl_tag,
    l_linestatus_o_valid             => PriceSummaryWriter_l_inst_l_linestatus_o_valid,
    l_linestatus_o_ready             => PriceSummaryWriter_l_inst_l_linestatus_o_ready,
    l_linestatus_o_dvalid            => PriceSummaryWriter_l_inst_l_linestatus_o_dvalid,
    l_linestatus_o_last              => PriceSummaryWriter_l_inst_l_linestatus_o_last,
    l_linestatus_o_length            => PriceSummaryWriter_l_inst_l_linestatus_o_length,
    l_linestatus_o_count             => PriceSummaryWriter_l_inst_l_linestatus_o_count,
    l_linestatus_o_chars_valid       => PriceSummaryWriter_l_inst_l_linestatus_o_chars_valid,
    l_linestatus_o_chars_ready       => PriceSummaryWriter_l_inst_l_linestatus_o_chars_ready,
    l_linestatus_o_chars_dvalid      => PriceSummaryWriter_l_inst_l_linestatus_o_chars_dvalid,
    l_linestatus_o_chars_last        => PriceSummaryWriter_l_inst_l_linestatus_o_chars_last,
    l_linestatus_o_chars             => PriceSummaryWriter_l_inst_l_linestatus_o_chars,
    l_linestatus_o_chars_count       => PriceSummaryWriter_l_inst_l_linestatus_o_chars_count,
    l_linestatus_o_bus_wreq_valid    => PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_valid,
    l_linestatus_o_bus_wreq_ready    => PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_ready,
    l_linestatus_o_bus_wreq_addr     => PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_addr,
    l_linestatus_o_bus_wreq_len      => PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_len,
    l_linestatus_o_bus_wdat_valid    => PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_valid,
    l_linestatus_o_bus_wdat_ready    => PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_ready,
    l_linestatus_o_bus_wdat_data     => PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_data,
    l_linestatus_o_bus_wdat_strobe   => PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_strobe,
    l_linestatus_o_bus_wdat_last     => PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_last,
    l_linestatus_o_cmd_valid         => PriceSummaryWriter_l_inst_l_linestatus_o_cmd_valid,
    l_linestatus_o_cmd_ready         => PriceSummaryWriter_l_inst_l_linestatus_o_cmd_ready,
    l_linestatus_o_cmd_firstIdx      => PriceSummaryWriter_l_inst_l_linestatus_o_cmd_firstIdx,
    l_linestatus_o_cmd_lastIdx       => PriceSummaryWriter_l_inst_l_linestatus_o_cmd_lastIdx,
    l_linestatus_o_cmd_ctrl          => PriceSummaryWriter_l_inst_l_linestatus_o_cmd_ctrl,
    l_linestatus_o_cmd_tag           => PriceSummaryWriter_l_inst_l_linestatus_o_cmd_tag,
    l_linestatus_o_unl_valid         => PriceSummaryWriter_l_inst_l_linestatus_o_unl_valid,
    l_linestatus_o_unl_ready         => PriceSummaryWriter_l_inst_l_linestatus_o_unl_ready,
    l_linestatus_o_unl_tag           => PriceSummaryWriter_l_inst_l_linestatus_o_unl_tag,
    l_sum_qty_valid                  => PriceSummaryWriter_l_inst_l_sum_qty_valid,
    l_sum_qty_ready                  => PriceSummaryWriter_l_inst_l_sum_qty_ready,
    l_sum_qty_dvalid                 => PriceSummaryWriter_l_inst_l_sum_qty_dvalid,
    l_sum_qty_last                   => PriceSummaryWriter_l_inst_l_sum_qty_last,
    l_sum_qty                        => PriceSummaryWriter_l_inst_l_sum_qty,
    l_sum_qty_bus_wreq_valid         => PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_valid,
    l_sum_qty_bus_wreq_ready         => PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_ready,
    l_sum_qty_bus_wreq_addr          => PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_addr,
    l_sum_qty_bus_wreq_len           => PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_len,
    l_sum_qty_bus_wdat_valid         => PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_valid,
    l_sum_qty_bus_wdat_ready         => PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_ready,
    l_sum_qty_bus_wdat_data          => PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_data,
    l_sum_qty_bus_wdat_strobe        => PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_strobe,
    l_sum_qty_bus_wdat_last          => PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_last,
    l_sum_qty_cmd_valid              => PriceSummaryWriter_l_inst_l_sum_qty_cmd_valid,
    l_sum_qty_cmd_ready              => PriceSummaryWriter_l_inst_l_sum_qty_cmd_ready,
    l_sum_qty_cmd_firstIdx           => PriceSummaryWriter_l_inst_l_sum_qty_cmd_firstIdx,
    l_sum_qty_cmd_lastIdx            => PriceSummaryWriter_l_inst_l_sum_qty_cmd_lastIdx,
    l_sum_qty_cmd_ctrl               => PriceSummaryWriter_l_inst_l_sum_qty_cmd_ctrl,
    l_sum_qty_cmd_tag                => PriceSummaryWriter_l_inst_l_sum_qty_cmd_tag,
    l_sum_qty_unl_valid              => PriceSummaryWriter_l_inst_l_sum_qty_unl_valid,
    l_sum_qty_unl_ready              => PriceSummaryWriter_l_inst_l_sum_qty_unl_ready,
    l_sum_qty_unl_tag                => PriceSummaryWriter_l_inst_l_sum_qty_unl_tag,
    l_sum_base_price_valid           => PriceSummaryWriter_l_inst_l_sum_base_price_valid,
    l_sum_base_price_ready           => PriceSummaryWriter_l_inst_l_sum_base_price_ready,
    l_sum_base_price_dvalid          => PriceSummaryWriter_l_inst_l_sum_base_price_dvalid,
    l_sum_base_price_last            => PriceSummaryWriter_l_inst_l_sum_base_price_last,
    l_sum_base_price                 => PriceSummaryWriter_l_inst_l_sum_base_price,
    l_sum_base_price_bus_wreq_valid  => PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_valid,
    l_sum_base_price_bus_wreq_ready  => PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_ready,
    l_sum_base_price_bus_wreq_addr   => PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_addr,
    l_sum_base_price_bus_wreq_len    => PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_len,
    l_sum_base_price_bus_wdat_valid  => PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_valid,
    l_sum_base_price_bus_wdat_ready  => PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_ready,
    l_sum_base_price_bus_wdat_data   => PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_data,
    l_sum_base_price_bus_wdat_strobe => PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_strobe,
    l_sum_base_price_bus_wdat_last   => PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_last,
    l_sum_base_price_cmd_valid       => PriceSummaryWriter_l_inst_l_sum_base_price_cmd_valid,
    l_sum_base_price_cmd_ready       => PriceSummaryWriter_l_inst_l_sum_base_price_cmd_ready,
    l_sum_base_price_cmd_firstIdx    => PriceSummaryWriter_l_inst_l_sum_base_price_cmd_firstIdx,
    l_sum_base_price_cmd_lastIdx     => PriceSummaryWriter_l_inst_l_sum_base_price_cmd_lastIdx,
    l_sum_base_price_cmd_ctrl        => PriceSummaryWriter_l_inst_l_sum_base_price_cmd_ctrl,
    l_sum_base_price_cmd_tag         => PriceSummaryWriter_l_inst_l_sum_base_price_cmd_tag,
    l_sum_base_price_unl_valid       => PriceSummaryWriter_l_inst_l_sum_base_price_unl_valid,
    l_sum_base_price_unl_ready       => PriceSummaryWriter_l_inst_l_sum_base_price_unl_ready,
    l_sum_base_price_unl_tag         => PriceSummaryWriter_l_inst_l_sum_base_price_unl_tag,
    l_sum_disc_price_valid           => PriceSummaryWriter_l_inst_l_sum_disc_price_valid,
    l_sum_disc_price_ready           => PriceSummaryWriter_l_inst_l_sum_disc_price_ready,
    l_sum_disc_price_dvalid          => PriceSummaryWriter_l_inst_l_sum_disc_price_dvalid,
    l_sum_disc_price_last            => PriceSummaryWriter_l_inst_l_sum_disc_price_last,
    l_sum_disc_price                 => PriceSummaryWriter_l_inst_l_sum_disc_price,
    l_sum_disc_price_bus_wreq_valid  => PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_valid,
    l_sum_disc_price_bus_wreq_ready  => PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_ready,
    l_sum_disc_price_bus_wreq_addr   => PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_addr,
    l_sum_disc_price_bus_wreq_len    => PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_len,
    l_sum_disc_price_bus_wdat_valid  => PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_valid,
    l_sum_disc_price_bus_wdat_ready  => PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_ready,
    l_sum_disc_price_bus_wdat_data   => PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_data,
    l_sum_disc_price_bus_wdat_strobe => PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_strobe,
    l_sum_disc_price_bus_wdat_last   => PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_last,
    l_sum_disc_price_cmd_valid       => PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_valid,
    l_sum_disc_price_cmd_ready       => PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_ready,
    l_sum_disc_price_cmd_firstIdx    => PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_firstIdx,
    l_sum_disc_price_cmd_lastIdx     => PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_lastIdx,
    l_sum_disc_price_cmd_ctrl        => PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_ctrl,
    l_sum_disc_price_cmd_tag         => PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_tag,
    l_sum_disc_price_unl_valid       => PriceSummaryWriter_l_inst_l_sum_disc_price_unl_valid,
    l_sum_disc_price_unl_ready       => PriceSummaryWriter_l_inst_l_sum_disc_price_unl_ready,
    l_sum_disc_price_unl_tag         => PriceSummaryWriter_l_inst_l_sum_disc_price_unl_tag,
    l_sum_charge_valid               => PriceSummaryWriter_l_inst_l_sum_charge_valid,
    l_sum_charge_ready               => PriceSummaryWriter_l_inst_l_sum_charge_ready,
    l_sum_charge_dvalid              => PriceSummaryWriter_l_inst_l_sum_charge_dvalid,
    l_sum_charge_last                => PriceSummaryWriter_l_inst_l_sum_charge_last,
    l_sum_charge                     => PriceSummaryWriter_l_inst_l_sum_charge,
    l_sum_charge_bus_wreq_valid      => PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_valid,
    l_sum_charge_bus_wreq_ready      => PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_ready,
    l_sum_charge_bus_wreq_addr       => PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_addr,
    l_sum_charge_bus_wreq_len        => PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_len,
    l_sum_charge_bus_wdat_valid      => PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_valid,
    l_sum_charge_bus_wdat_ready      => PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_ready,
    l_sum_charge_bus_wdat_data       => PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_data,
    l_sum_charge_bus_wdat_strobe     => PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_strobe,
    l_sum_charge_bus_wdat_last       => PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_last,
    l_sum_charge_cmd_valid           => PriceSummaryWriter_l_inst_l_sum_charge_cmd_valid,
    l_sum_charge_cmd_ready           => PriceSummaryWriter_l_inst_l_sum_charge_cmd_ready,
    l_sum_charge_cmd_firstIdx        => PriceSummaryWriter_l_inst_l_sum_charge_cmd_firstIdx,
    l_sum_charge_cmd_lastIdx         => PriceSummaryWriter_l_inst_l_sum_charge_cmd_lastIdx,
    l_sum_charge_cmd_ctrl            => PriceSummaryWriter_l_inst_l_sum_charge_cmd_ctrl,
    l_sum_charge_cmd_tag             => PriceSummaryWriter_l_inst_l_sum_charge_cmd_tag,
    l_sum_charge_unl_valid           => PriceSummaryWriter_l_inst_l_sum_charge_unl_valid,
    l_sum_charge_unl_ready           => PriceSummaryWriter_l_inst_l_sum_charge_unl_ready,
    l_sum_charge_unl_tag             => PriceSummaryWriter_l_inst_l_sum_charge_unl_tag,
    l_avg_qty_valid                  => PriceSummaryWriter_l_inst_l_avg_qty_valid,
    l_avg_qty_ready                  => PriceSummaryWriter_l_inst_l_avg_qty_ready,
    l_avg_qty_dvalid                 => PriceSummaryWriter_l_inst_l_avg_qty_dvalid,
    l_avg_qty_last                   => PriceSummaryWriter_l_inst_l_avg_qty_last,
    l_avg_qty                        => PriceSummaryWriter_l_inst_l_avg_qty,
    l_avg_qty_bus_wreq_valid         => PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_valid,
    l_avg_qty_bus_wreq_ready         => PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_ready,
    l_avg_qty_bus_wreq_addr          => PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_addr,
    l_avg_qty_bus_wreq_len           => PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_len,
    l_avg_qty_bus_wdat_valid         => PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_valid,
    l_avg_qty_bus_wdat_ready         => PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_ready,
    l_avg_qty_bus_wdat_data          => PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_data,
    l_avg_qty_bus_wdat_strobe        => PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_strobe,
    l_avg_qty_bus_wdat_last          => PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_last,
    l_avg_qty_cmd_valid              => PriceSummaryWriter_l_inst_l_avg_qty_cmd_valid,
    l_avg_qty_cmd_ready              => PriceSummaryWriter_l_inst_l_avg_qty_cmd_ready,
    l_avg_qty_cmd_firstIdx           => PriceSummaryWriter_l_inst_l_avg_qty_cmd_firstIdx,
    l_avg_qty_cmd_lastIdx            => PriceSummaryWriter_l_inst_l_avg_qty_cmd_lastIdx,
    l_avg_qty_cmd_ctrl               => PriceSummaryWriter_l_inst_l_avg_qty_cmd_ctrl,
    l_avg_qty_cmd_tag                => PriceSummaryWriter_l_inst_l_avg_qty_cmd_tag,
    l_avg_qty_unl_valid              => PriceSummaryWriter_l_inst_l_avg_qty_unl_valid,
    l_avg_qty_unl_ready              => PriceSummaryWriter_l_inst_l_avg_qty_unl_ready,
    l_avg_qty_unl_tag                => PriceSummaryWriter_l_inst_l_avg_qty_unl_tag,
    l_avg_price_valid                => PriceSummaryWriter_l_inst_l_avg_price_valid,
    l_avg_price_ready                => PriceSummaryWriter_l_inst_l_avg_price_ready,
    l_avg_price_dvalid               => PriceSummaryWriter_l_inst_l_avg_price_dvalid,
    l_avg_price_last                 => PriceSummaryWriter_l_inst_l_avg_price_last,
    l_avg_price                      => PriceSummaryWriter_l_inst_l_avg_price,
    l_avg_price_bus_wreq_valid       => PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_valid,
    l_avg_price_bus_wreq_ready       => PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_ready,
    l_avg_price_bus_wreq_addr        => PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_addr,
    l_avg_price_bus_wreq_len         => PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_len,
    l_avg_price_bus_wdat_valid       => PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_valid,
    l_avg_price_bus_wdat_ready       => PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_ready,
    l_avg_price_bus_wdat_data        => PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_data,
    l_avg_price_bus_wdat_strobe      => PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_strobe,
    l_avg_price_bus_wdat_last        => PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_last,
    l_avg_price_cmd_valid            => PriceSummaryWriter_l_inst_l_avg_price_cmd_valid,
    l_avg_price_cmd_ready            => PriceSummaryWriter_l_inst_l_avg_price_cmd_ready,
    l_avg_price_cmd_firstIdx         => PriceSummaryWriter_l_inst_l_avg_price_cmd_firstIdx,
    l_avg_price_cmd_lastIdx          => PriceSummaryWriter_l_inst_l_avg_price_cmd_lastIdx,
    l_avg_price_cmd_ctrl             => PriceSummaryWriter_l_inst_l_avg_price_cmd_ctrl,
    l_avg_price_cmd_tag              => PriceSummaryWriter_l_inst_l_avg_price_cmd_tag,
    l_avg_price_unl_valid            => PriceSummaryWriter_l_inst_l_avg_price_unl_valid,
    l_avg_price_unl_ready            => PriceSummaryWriter_l_inst_l_avg_price_unl_ready,
    l_avg_price_unl_tag              => PriceSummaryWriter_l_inst_l_avg_price_unl_tag,
    l_avg_disc_valid                 => PriceSummaryWriter_l_inst_l_avg_disc_valid,
    l_avg_disc_ready                 => PriceSummaryWriter_l_inst_l_avg_disc_ready,
    l_avg_disc_dvalid                => PriceSummaryWriter_l_inst_l_avg_disc_dvalid,
    l_avg_disc_last                  => PriceSummaryWriter_l_inst_l_avg_disc_last,
    l_avg_disc                       => PriceSummaryWriter_l_inst_l_avg_disc,
    l_avg_disc_bus_wreq_valid        => PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_valid,
    l_avg_disc_bus_wreq_ready        => PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_ready,
    l_avg_disc_bus_wreq_addr         => PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_addr,
    l_avg_disc_bus_wreq_len          => PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_len,
    l_avg_disc_bus_wdat_valid        => PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_valid,
    l_avg_disc_bus_wdat_ready        => PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_ready,
    l_avg_disc_bus_wdat_data         => PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_data,
    l_avg_disc_bus_wdat_strobe       => PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_strobe,
    l_avg_disc_bus_wdat_last         => PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_last,
    l_avg_disc_cmd_valid             => PriceSummaryWriter_l_inst_l_avg_disc_cmd_valid,
    l_avg_disc_cmd_ready             => PriceSummaryWriter_l_inst_l_avg_disc_cmd_ready,
    l_avg_disc_cmd_firstIdx          => PriceSummaryWriter_l_inst_l_avg_disc_cmd_firstIdx,
    l_avg_disc_cmd_lastIdx           => PriceSummaryWriter_l_inst_l_avg_disc_cmd_lastIdx,
    l_avg_disc_cmd_ctrl              => PriceSummaryWriter_l_inst_l_avg_disc_cmd_ctrl,
    l_avg_disc_cmd_tag               => PriceSummaryWriter_l_inst_l_avg_disc_cmd_tag,
    l_avg_disc_unl_valid             => PriceSummaryWriter_l_inst_l_avg_disc_unl_valid,
    l_avg_disc_unl_ready             => PriceSummaryWriter_l_inst_l_avg_disc_unl_ready,
    l_avg_disc_unl_tag               => PriceSummaryWriter_l_inst_l_avg_disc_unl_tag,
    l_count_order_valid              => PriceSummaryWriter_l_inst_l_count_order_valid,
    l_count_order_ready              => PriceSummaryWriter_l_inst_l_count_order_ready,
    l_count_order_dvalid             => PriceSummaryWriter_l_inst_l_count_order_dvalid,
    l_count_order_last               => PriceSummaryWriter_l_inst_l_count_order_last,
    l_count_order                    => PriceSummaryWriter_l_inst_l_count_order,
    l_count_order_bus_wreq_valid     => PriceSummaryWriter_l_inst_l_count_order_bus_wreq_valid,
    l_count_order_bus_wreq_ready     => PriceSummaryWriter_l_inst_l_count_order_bus_wreq_ready,
    l_count_order_bus_wreq_addr      => PriceSummaryWriter_l_inst_l_count_order_bus_wreq_addr,
    l_count_order_bus_wreq_len       => PriceSummaryWriter_l_inst_l_count_order_bus_wreq_len,
    l_count_order_bus_wdat_valid     => PriceSummaryWriter_l_inst_l_count_order_bus_wdat_valid,
    l_count_order_bus_wdat_ready     => PriceSummaryWriter_l_inst_l_count_order_bus_wdat_ready,
    l_count_order_bus_wdat_data      => PriceSummaryWriter_l_inst_l_count_order_bus_wdat_data,
    l_count_order_bus_wdat_strobe    => PriceSummaryWriter_l_inst_l_count_order_bus_wdat_strobe,
    l_count_order_bus_wdat_last      => PriceSummaryWriter_l_inst_l_count_order_bus_wdat_last,
    l_count_order_cmd_valid          => PriceSummaryWriter_l_inst_l_count_order_cmd_valid,
    l_count_order_cmd_ready          => PriceSummaryWriter_l_inst_l_count_order_cmd_ready,
    l_count_order_cmd_firstIdx       => PriceSummaryWriter_l_inst_l_count_order_cmd_firstIdx,
    l_count_order_cmd_lastIdx        => PriceSummaryWriter_l_inst_l_count_order_cmd_lastIdx,
    l_count_order_cmd_ctrl           => PriceSummaryWriter_l_inst_l_count_order_cmd_ctrl,
    l_count_order_cmd_tag            => PriceSummaryWriter_l_inst_l_count_order_cmd_tag,
    l_count_order_unl_valid          => PriceSummaryWriter_l_inst_l_count_order_unl_valid,
    l_count_order_unl_ready          => PriceSummaryWriter_l_inst_l_count_order_unl_ready,
    l_count_order_unl_tag            => PriceSummaryWriter_l_inst_l_count_order_unl_tag
  );

  WRAW64DW512LW8BS1BM16_inst : BusWriteArbiterVec
  generic map(
    BUS_ADDR_WIDTH  => BUS_ADDR_WIDTH,
    BUS_DATA_WIDTH  => BUS_DATA_WIDTH,
    BUS_LEN_WIDTH   => BUS_LEN_WIDTH,
    NUM_SLAVE_PORTS => 10,
    ARB_METHOD      => "RR-STICKY",
    MAX_OUTSTANDING => 4,
    RAM_CONFIG      => "",
    SLV_REQ_SLICES  => true,
    MST_REQ_SLICE   => true,
    MST_DAT_SLICE   => true,
    SLV_DAT_SLICES  => true
  )
  port map(
    bcd_clk         => bcd_clk,
    bcd_reset       => bcd_reset,
    mst_wreq_valid  => WRAW64DW512LW8BS1BM16_inst_mst_wreq_valid,
    mst_wreq_ready  => WRAW64DW512LW8BS1BM16_inst_mst_wreq_ready,
    mst_wreq_addr   => WRAW64DW512LW8BS1BM16_inst_mst_wreq_addr,
    mst_wreq_len    => WRAW64DW512LW8BS1BM16_inst_mst_wreq_len,
    mst_wdat_valid  => WRAW64DW512LW8BS1BM16_inst_mst_wdat_valid,
    mst_wdat_ready  => WRAW64DW512LW8BS1BM16_inst_mst_wdat_ready,
    mst_wdat_data   => WRAW64DW512LW8BS1BM16_inst_mst_wdat_data,
    mst_wdat_strobe => WRAW64DW512LW8BS1BM16_inst_mst_wdat_strobe,
    mst_wdat_last   => WRAW64DW512LW8BS1BM16_inst_mst_wdat_last,
    bsv_wreq_valid  => WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid,
    bsv_wreq_ready  => WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready,
    bsv_wreq_len    => WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len,
    bsv_wreq_addr   => WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr,
    bsv_wdat_valid  => WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid,
    bsv_wdat_strobe => WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe,
    bsv_wdat_ready  => WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready,
    bsv_wdat_last   => WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last,
    bsv_wdat_data   => WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data
  );

  wr_mst_wreq_valid                                                                                                   <= WRAW64DW512LW8BS1BM16_inst_mst_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_mst_wreq_ready                                                                           <= wr_mst_wreq_ready;
  wr_mst_wreq_addr                                                                                                    <= WRAW64DW512LW8BS1BM16_inst_mst_wreq_addr;
  wr_mst_wreq_len                                                                                                     <= WRAW64DW512LW8BS1BM16_inst_mst_wreq_len;
  wr_mst_wdat_valid                                                                                                   <= WRAW64DW512LW8BS1BM16_inst_mst_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_mst_wdat_ready                                                                           <= wr_mst_wdat_ready;
  wr_mst_wdat_data                                                                                                    <= WRAW64DW512LW8BS1BM16_inst_mst_wdat_data;
  wr_mst_wdat_strobe                                                                                                  <= WRAW64DW512LW8BS1BM16_inst_mst_wdat_strobe;
  wr_mst_wdat_last                                                                                                    <= WRAW64DW512LW8BS1BM16_inst_mst_wdat_last;

  PriceSummaryWriter_Nucleus_inst_l_returnflag_o_unl_valid                                                            <= PriceSummaryWriter_l_inst_l_returnflag_o_unl_valid;
  PriceSummaryWriter_l_inst_l_returnflag_o_unl_ready                                                                  <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_unl_ready;
  PriceSummaryWriter_Nucleus_inst_l_returnflag_o_unl_tag                                                              <= PriceSummaryWriter_l_inst_l_returnflag_o_unl_tag;

  PriceSummaryWriter_Nucleus_inst_l_linestatus_o_unl_valid                                                            <= PriceSummaryWriter_l_inst_l_linestatus_o_unl_valid;
  PriceSummaryWriter_l_inst_l_linestatus_o_unl_ready                                                                  <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_unl_ready;
  PriceSummaryWriter_Nucleus_inst_l_linestatus_o_unl_tag                                                              <= PriceSummaryWriter_l_inst_l_linestatus_o_unl_tag;

  PriceSummaryWriter_Nucleus_inst_l_sum_qty_unl_valid                                                                 <= PriceSummaryWriter_l_inst_l_sum_qty_unl_valid;
  PriceSummaryWriter_l_inst_l_sum_qty_unl_ready                                                                       <= PriceSummaryWriter_Nucleus_inst_l_sum_qty_unl_ready;
  PriceSummaryWriter_Nucleus_inst_l_sum_qty_unl_tag                                                                   <= PriceSummaryWriter_l_inst_l_sum_qty_unl_tag;

  PriceSummaryWriter_Nucleus_inst_l_sum_base_price_unl_valid                                                          <= PriceSummaryWriter_l_inst_l_sum_base_price_unl_valid;
  PriceSummaryWriter_l_inst_l_sum_base_price_unl_ready                                                                <= PriceSummaryWriter_Nucleus_inst_l_sum_base_price_unl_ready;
  PriceSummaryWriter_Nucleus_inst_l_sum_base_price_unl_tag                                                            <= PriceSummaryWriter_l_inst_l_sum_base_price_unl_tag;

  PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_unl_valid                                                          <= PriceSummaryWriter_l_inst_l_sum_disc_price_unl_valid;
  PriceSummaryWriter_l_inst_l_sum_disc_price_unl_ready                                                                <= PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_unl_ready;
  PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_unl_tag                                                            <= PriceSummaryWriter_l_inst_l_sum_disc_price_unl_tag;

  PriceSummaryWriter_Nucleus_inst_l_sum_charge_unl_valid                                                              <= PriceSummaryWriter_l_inst_l_sum_charge_unl_valid;
  PriceSummaryWriter_l_inst_l_sum_charge_unl_ready                                                                    <= PriceSummaryWriter_Nucleus_inst_l_sum_charge_unl_ready;
  PriceSummaryWriter_Nucleus_inst_l_sum_charge_unl_tag                                                                <= PriceSummaryWriter_l_inst_l_sum_charge_unl_tag;

  PriceSummaryWriter_Nucleus_inst_l_avg_qty_unl_valid                                                                 <= PriceSummaryWriter_l_inst_l_avg_qty_unl_valid;
  PriceSummaryWriter_l_inst_l_avg_qty_unl_ready                                                                       <= PriceSummaryWriter_Nucleus_inst_l_avg_qty_unl_ready;
  PriceSummaryWriter_Nucleus_inst_l_avg_qty_unl_tag                                                                   <= PriceSummaryWriter_l_inst_l_avg_qty_unl_tag;

  PriceSummaryWriter_Nucleus_inst_l_avg_price_unl_valid                                                               <= PriceSummaryWriter_l_inst_l_avg_price_unl_valid;
  PriceSummaryWriter_l_inst_l_avg_price_unl_ready                                                                     <= PriceSummaryWriter_Nucleus_inst_l_avg_price_unl_ready;
  PriceSummaryWriter_Nucleus_inst_l_avg_price_unl_tag                                                                 <= PriceSummaryWriter_l_inst_l_avg_price_unl_tag;

  PriceSummaryWriter_Nucleus_inst_l_avg_disc_unl_valid                                                                <= PriceSummaryWriter_l_inst_l_avg_disc_unl_valid;
  PriceSummaryWriter_l_inst_l_avg_disc_unl_ready                                                                      <= PriceSummaryWriter_Nucleus_inst_l_avg_disc_unl_ready;
  PriceSummaryWriter_Nucleus_inst_l_avg_disc_unl_tag                                                                  <= PriceSummaryWriter_l_inst_l_avg_disc_unl_tag;

  PriceSummaryWriter_Nucleus_inst_l_count_order_unl_valid                                                             <= PriceSummaryWriter_l_inst_l_count_order_unl_valid;
  PriceSummaryWriter_l_inst_l_count_order_unl_ready                                                                   <= PriceSummaryWriter_Nucleus_inst_l_count_order_unl_ready;
  PriceSummaryWriter_Nucleus_inst_l_count_order_unl_tag                                                               <= PriceSummaryWriter_l_inst_l_count_order_unl_tag;

  PriceSummaryWriter_l_inst_l_returnflag_o_valid                                                                      <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_valid;
  PriceSummaryWriter_Nucleus_inst_l_returnflag_o_ready                                                                <= PriceSummaryWriter_l_inst_l_returnflag_o_ready;
  PriceSummaryWriter_l_inst_l_returnflag_o_dvalid                                                                     <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_dvalid;
  PriceSummaryWriter_l_inst_l_returnflag_o_last                                                                       <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_last;
  PriceSummaryWriter_l_inst_l_returnflag_o_length                                                                     <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_length;
  PriceSummaryWriter_l_inst_l_returnflag_o_count                                                                      <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_count;
  PriceSummaryWriter_l_inst_l_returnflag_o_chars_valid                                                                <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_valid;
  PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_ready                                                          <= PriceSummaryWriter_l_inst_l_returnflag_o_chars_ready;
  PriceSummaryWriter_l_inst_l_returnflag_o_chars_dvalid                                                               <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_dvalid;
  PriceSummaryWriter_l_inst_l_returnflag_o_chars_last                                                                 <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_last;
  PriceSummaryWriter_l_inst_l_returnflag_o_chars                                                                      <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars;
  PriceSummaryWriter_l_inst_l_returnflag_o_chars_count                                                                <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_count;

  PriceSummaryWriter_l_inst_l_returnflag_o_cmd_valid                                                                  <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_valid;
  PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_ready                                                            <= PriceSummaryWriter_l_inst_l_returnflag_o_cmd_ready;
  PriceSummaryWriter_l_inst_l_returnflag_o_cmd_firstIdx                                                               <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_firstIdx;
  PriceSummaryWriter_l_inst_l_returnflag_o_cmd_lastIdx                                                                <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_lastIdx;
  PriceSummaryWriter_l_inst_l_returnflag_o_cmd_ctrl                                                                   <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_ctrl;
  PriceSummaryWriter_l_inst_l_returnflag_o_cmd_tag                                                                    <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_tag;

  PriceSummaryWriter_l_inst_l_linestatus_o_valid                                                                      <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_valid;
  PriceSummaryWriter_Nucleus_inst_l_linestatus_o_ready                                                                <= PriceSummaryWriter_l_inst_l_linestatus_o_ready;
  PriceSummaryWriter_l_inst_l_linestatus_o_dvalid                                                                     <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_dvalid;
  PriceSummaryWriter_l_inst_l_linestatus_o_last                                                                       <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_last;
  PriceSummaryWriter_l_inst_l_linestatus_o_length                                                                     <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_length;
  PriceSummaryWriter_l_inst_l_linestatus_o_count                                                                      <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_count;
  PriceSummaryWriter_l_inst_l_linestatus_o_chars_valid                                                                <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_valid;
  PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_ready                                                          <= PriceSummaryWriter_l_inst_l_linestatus_o_chars_ready;
  PriceSummaryWriter_l_inst_l_linestatus_o_chars_dvalid                                                               <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_dvalid;
  PriceSummaryWriter_l_inst_l_linestatus_o_chars_last                                                                 <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_last;
  PriceSummaryWriter_l_inst_l_linestatus_o_chars                                                                      <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars;
  PriceSummaryWriter_l_inst_l_linestatus_o_chars_count                                                                <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_count;

  PriceSummaryWriter_l_inst_l_linestatus_o_cmd_valid                                                                  <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_valid;
  PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_ready                                                            <= PriceSummaryWriter_l_inst_l_linestatus_o_cmd_ready;
  PriceSummaryWriter_l_inst_l_linestatus_o_cmd_firstIdx                                                               <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_firstIdx;
  PriceSummaryWriter_l_inst_l_linestatus_o_cmd_lastIdx                                                                <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_lastIdx;
  PriceSummaryWriter_l_inst_l_linestatus_o_cmd_ctrl                                                                   <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_ctrl;
  PriceSummaryWriter_l_inst_l_linestatus_o_cmd_tag                                                                    <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_tag;

  PriceSummaryWriter_l_inst_l_sum_qty_valid                                                                           <= PriceSummaryWriter_Nucleus_inst_l_sum_qty_valid;
  PriceSummaryWriter_Nucleus_inst_l_sum_qty_ready                                                                     <= PriceSummaryWriter_l_inst_l_sum_qty_ready;
  PriceSummaryWriter_l_inst_l_sum_qty_dvalid                                                                          <= PriceSummaryWriter_Nucleus_inst_l_sum_qty_dvalid;
  PriceSummaryWriter_l_inst_l_sum_qty_last                                                                            <= PriceSummaryWriter_Nucleus_inst_l_sum_qty_last;
  PriceSummaryWriter_l_inst_l_sum_qty                                                                                 <= PriceSummaryWriter_Nucleus_inst_l_sum_qty;

  PriceSummaryWriter_l_inst_l_sum_qty_cmd_valid                                                                       <= PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_valid;
  PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_ready                                                                 <= PriceSummaryWriter_l_inst_l_sum_qty_cmd_ready;
  PriceSummaryWriter_l_inst_l_sum_qty_cmd_firstIdx                                                                    <= PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_firstIdx;
  PriceSummaryWriter_l_inst_l_sum_qty_cmd_lastIdx                                                                     <= PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_lastIdx;
  PriceSummaryWriter_l_inst_l_sum_qty_cmd_ctrl                                                                        <= PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_ctrl;
  PriceSummaryWriter_l_inst_l_sum_qty_cmd_tag                                                                         <= PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_tag;

  PriceSummaryWriter_l_inst_l_sum_base_price_valid                                                                    <= PriceSummaryWriter_Nucleus_inst_l_sum_base_price_valid;
  PriceSummaryWriter_Nucleus_inst_l_sum_base_price_ready                                                              <= PriceSummaryWriter_l_inst_l_sum_base_price_ready;
  PriceSummaryWriter_l_inst_l_sum_base_price_dvalid                                                                   <= PriceSummaryWriter_Nucleus_inst_l_sum_base_price_dvalid;
  PriceSummaryWriter_l_inst_l_sum_base_price_last                                                                     <= PriceSummaryWriter_Nucleus_inst_l_sum_base_price_last;
  PriceSummaryWriter_l_inst_l_sum_base_price                                                                          <= PriceSummaryWriter_Nucleus_inst_l_sum_base_price;

  PriceSummaryWriter_l_inst_l_sum_base_price_cmd_valid                                                                <= PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_valid;
  PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_ready                                                          <= PriceSummaryWriter_l_inst_l_sum_base_price_cmd_ready;
  PriceSummaryWriter_l_inst_l_sum_base_price_cmd_firstIdx                                                             <= PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_firstIdx;
  PriceSummaryWriter_l_inst_l_sum_base_price_cmd_lastIdx                                                              <= PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_lastIdx;
  PriceSummaryWriter_l_inst_l_sum_base_price_cmd_ctrl                                                                 <= PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_ctrl;
  PriceSummaryWriter_l_inst_l_sum_base_price_cmd_tag                                                                  <= PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_tag;

  PriceSummaryWriter_l_inst_l_sum_disc_price_valid                                                                    <= PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_valid;
  PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_ready                                                              <= PriceSummaryWriter_l_inst_l_sum_disc_price_ready;
  PriceSummaryWriter_l_inst_l_sum_disc_price_dvalid                                                                   <= PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_dvalid;
  PriceSummaryWriter_l_inst_l_sum_disc_price_last                                                                     <= PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_last;
  PriceSummaryWriter_l_inst_l_sum_disc_price                                                                          <= PriceSummaryWriter_Nucleus_inst_l_sum_disc_price;

  PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_valid                                                                <= PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_valid;
  PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_ready                                                          <= PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_ready;
  PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_firstIdx                                                             <= PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_firstIdx;
  PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_lastIdx                                                              <= PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_lastIdx;
  PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_ctrl                                                                 <= PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_ctrl;
  PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_tag                                                                  <= PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_tag;

  PriceSummaryWriter_l_inst_l_sum_charge_valid                                                                        <= PriceSummaryWriter_Nucleus_inst_l_sum_charge_valid;
  PriceSummaryWriter_Nucleus_inst_l_sum_charge_ready                                                                  <= PriceSummaryWriter_l_inst_l_sum_charge_ready;
  PriceSummaryWriter_l_inst_l_sum_charge_dvalid                                                                       <= PriceSummaryWriter_Nucleus_inst_l_sum_charge_dvalid;
  PriceSummaryWriter_l_inst_l_sum_charge_last                                                                         <= PriceSummaryWriter_Nucleus_inst_l_sum_charge_last;
  PriceSummaryWriter_l_inst_l_sum_charge                                                                              <= PriceSummaryWriter_Nucleus_inst_l_sum_charge;

  PriceSummaryWriter_l_inst_l_sum_charge_cmd_valid                                                                    <= PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_valid;
  PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_ready                                                              <= PriceSummaryWriter_l_inst_l_sum_charge_cmd_ready;
  PriceSummaryWriter_l_inst_l_sum_charge_cmd_firstIdx                                                                 <= PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_firstIdx;
  PriceSummaryWriter_l_inst_l_sum_charge_cmd_lastIdx                                                                  <= PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_lastIdx;
  PriceSummaryWriter_l_inst_l_sum_charge_cmd_ctrl                                                                     <= PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_ctrl;
  PriceSummaryWriter_l_inst_l_sum_charge_cmd_tag                                                                      <= PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_tag;

  PriceSummaryWriter_l_inst_l_avg_qty_valid                                                                           <= PriceSummaryWriter_Nucleus_inst_l_avg_qty_valid;
  PriceSummaryWriter_Nucleus_inst_l_avg_qty_ready                                                                     <= PriceSummaryWriter_l_inst_l_avg_qty_ready;
  PriceSummaryWriter_l_inst_l_avg_qty_dvalid                                                                          <= PriceSummaryWriter_Nucleus_inst_l_avg_qty_dvalid;
  PriceSummaryWriter_l_inst_l_avg_qty_last                                                                            <= PriceSummaryWriter_Nucleus_inst_l_avg_qty_last;
  PriceSummaryWriter_l_inst_l_avg_qty                                                                                 <= PriceSummaryWriter_Nucleus_inst_l_avg_qty;

  PriceSummaryWriter_l_inst_l_avg_qty_cmd_valid                                                                       <= PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_valid;
  PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_ready                                                                 <= PriceSummaryWriter_l_inst_l_avg_qty_cmd_ready;
  PriceSummaryWriter_l_inst_l_avg_qty_cmd_firstIdx                                                                    <= PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_firstIdx;
  PriceSummaryWriter_l_inst_l_avg_qty_cmd_lastIdx                                                                     <= PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_lastIdx;
  PriceSummaryWriter_l_inst_l_avg_qty_cmd_ctrl                                                                        <= PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_ctrl;
  PriceSummaryWriter_l_inst_l_avg_qty_cmd_tag                                                                         <= PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_tag;

  PriceSummaryWriter_l_inst_l_avg_price_valid                                                                         <= PriceSummaryWriter_Nucleus_inst_l_avg_price_valid;
  PriceSummaryWriter_Nucleus_inst_l_avg_price_ready                                                                   <= PriceSummaryWriter_l_inst_l_avg_price_ready;
  PriceSummaryWriter_l_inst_l_avg_price_dvalid                                                                        <= PriceSummaryWriter_Nucleus_inst_l_avg_price_dvalid;
  PriceSummaryWriter_l_inst_l_avg_price_last                                                                          <= PriceSummaryWriter_Nucleus_inst_l_avg_price_last;
  PriceSummaryWriter_l_inst_l_avg_price                                                                               <= PriceSummaryWriter_Nucleus_inst_l_avg_price;

  PriceSummaryWriter_l_inst_l_avg_price_cmd_valid                                                                     <= PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_valid;
  PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_ready                                                               <= PriceSummaryWriter_l_inst_l_avg_price_cmd_ready;
  PriceSummaryWriter_l_inst_l_avg_price_cmd_firstIdx                                                                  <= PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_firstIdx;
  PriceSummaryWriter_l_inst_l_avg_price_cmd_lastIdx                                                                   <= PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_lastIdx;
  PriceSummaryWriter_l_inst_l_avg_price_cmd_ctrl                                                                      <= PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_ctrl;
  PriceSummaryWriter_l_inst_l_avg_price_cmd_tag                                                                       <= PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_tag;

  PriceSummaryWriter_l_inst_l_avg_disc_valid                                                                          <= PriceSummaryWriter_Nucleus_inst_l_avg_disc_valid;
  PriceSummaryWriter_Nucleus_inst_l_avg_disc_ready                                                                    <= PriceSummaryWriter_l_inst_l_avg_disc_ready;
  PriceSummaryWriter_l_inst_l_avg_disc_dvalid                                                                         <= PriceSummaryWriter_Nucleus_inst_l_avg_disc_dvalid;
  PriceSummaryWriter_l_inst_l_avg_disc_last                                                                           <= PriceSummaryWriter_Nucleus_inst_l_avg_disc_last;
  PriceSummaryWriter_l_inst_l_avg_disc                                                                                <= PriceSummaryWriter_Nucleus_inst_l_avg_disc;

  PriceSummaryWriter_l_inst_l_avg_disc_cmd_valid                                                                      <= PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_valid;
  PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_ready                                                                <= PriceSummaryWriter_l_inst_l_avg_disc_cmd_ready;
  PriceSummaryWriter_l_inst_l_avg_disc_cmd_firstIdx                                                                   <= PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_firstIdx;
  PriceSummaryWriter_l_inst_l_avg_disc_cmd_lastIdx                                                                    <= PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_lastIdx;
  PriceSummaryWriter_l_inst_l_avg_disc_cmd_ctrl                                                                       <= PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_ctrl;
  PriceSummaryWriter_l_inst_l_avg_disc_cmd_tag                                                                        <= PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_tag;

  PriceSummaryWriter_l_inst_l_count_order_valid                                                                       <= PriceSummaryWriter_Nucleus_inst_l_count_order_valid;
  PriceSummaryWriter_Nucleus_inst_l_count_order_ready                                                                 <= PriceSummaryWriter_l_inst_l_count_order_ready;
  PriceSummaryWriter_l_inst_l_count_order_dvalid                                                                      <= PriceSummaryWriter_Nucleus_inst_l_count_order_dvalid;
  PriceSummaryWriter_l_inst_l_count_order_last                                                                        <= PriceSummaryWriter_Nucleus_inst_l_count_order_last;
  PriceSummaryWriter_l_inst_l_count_order                                                                             <= PriceSummaryWriter_Nucleus_inst_l_count_order;

  PriceSummaryWriter_l_inst_l_count_order_cmd_valid                                                                   <= PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_valid;
  PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_ready                                                             <= PriceSummaryWriter_l_inst_l_count_order_cmd_ready;
  PriceSummaryWriter_l_inst_l_count_order_cmd_firstIdx                                                                <= PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_firstIdx;
  PriceSummaryWriter_l_inst_l_count_order_cmd_lastIdx                                                                 <= PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_lastIdx;
  PriceSummaryWriter_l_inst_l_count_order_cmd_ctrl                                                                    <= PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_ctrl;
  PriceSummaryWriter_l_inst_l_count_order_cmd_tag                                                                     <= PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_tag;

  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid(0)                                                                        <= PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid(1)                                                                        <= PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid(2)                                                                        <= PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid(3)                                                                        <= PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid(4)                                                                        <= PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid(5)                                                                        <= PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid(6)                                                                        <= PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid(7)                                                                        <= PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid(8)                                                                        <= PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid(9)                                                                        <= PriceSummaryWriter_l_inst_l_count_order_bus_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len(BUS_LEN_WIDTH - 1 downto 0)                                                 <= PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_len;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len(BUS_LEN_WIDTH + BUS_LEN_WIDTH - 1 downto BUS_LEN_WIDTH)                     <= PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_len;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len(BUS_LEN_WIDTH * 2 + BUS_LEN_WIDTH - 1 downto BUS_LEN_WIDTH * 2)             <= PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_len;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len(BUS_LEN_WIDTH * 3 + BUS_LEN_WIDTH - 1 downto BUS_LEN_WIDTH * 3)             <= PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_len;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len(BUS_LEN_WIDTH * 4 + BUS_LEN_WIDTH - 1 downto BUS_LEN_WIDTH * 4)             <= PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_len;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len(BUS_LEN_WIDTH * 5 + BUS_LEN_WIDTH - 1 downto BUS_LEN_WIDTH * 5)             <= PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_len;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len(BUS_LEN_WIDTH * 6 + BUS_LEN_WIDTH - 1 downto BUS_LEN_WIDTH * 6)             <= PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_len;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len(BUS_LEN_WIDTH * 7 + BUS_LEN_WIDTH - 1 downto BUS_LEN_WIDTH * 7)             <= PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_len;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len(BUS_LEN_WIDTH * 8 + BUS_LEN_WIDTH - 1 downto BUS_LEN_WIDTH * 8)             <= PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_len;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len(BUS_LEN_WIDTH * 9 + BUS_LEN_WIDTH - 1 downto BUS_LEN_WIDTH * 9)             <= PriceSummaryWriter_l_inst_l_count_order_bus_wreq_len;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr(BUS_ADDR_WIDTH - 1 downto 0)                                               <= PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_addr;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr(BUS_ADDR_WIDTH + BUS_ADDR_WIDTH - 1 downto BUS_ADDR_WIDTH)                 <= PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_addr;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr(BUS_ADDR_WIDTH * 2 + BUS_ADDR_WIDTH - 1 downto BUS_ADDR_WIDTH * 2)         <= PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_addr;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr(BUS_ADDR_WIDTH * 3 + BUS_ADDR_WIDTH - 1 downto BUS_ADDR_WIDTH * 3)         <= PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_addr;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr(BUS_ADDR_WIDTH * 4 + BUS_ADDR_WIDTH - 1 downto BUS_ADDR_WIDTH * 4)         <= PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_addr;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr(BUS_ADDR_WIDTH * 5 + BUS_ADDR_WIDTH - 1 downto BUS_ADDR_WIDTH * 5)         <= PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_addr;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr(BUS_ADDR_WIDTH * 6 + BUS_ADDR_WIDTH - 1 downto BUS_ADDR_WIDTH * 6)         <= PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_addr;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr(BUS_ADDR_WIDTH * 7 + BUS_ADDR_WIDTH - 1 downto BUS_ADDR_WIDTH * 7)         <= PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_addr;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr(BUS_ADDR_WIDTH * 8 + BUS_ADDR_WIDTH - 1 downto BUS_ADDR_WIDTH * 8)         <= PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_addr;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr(BUS_ADDR_WIDTH * 9 + BUS_ADDR_WIDTH - 1 downto BUS_ADDR_WIDTH * 9)         <= PriceSummaryWriter_l_inst_l_count_order_bus_wreq_addr;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid(0)                                                                        <= PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid(1)                                                                        <= PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid(2)                                                                        <= PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid(3)                                                                        <= PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid(4)                                                                        <= PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid(5)                                                                        <= PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid(6)                                                                        <= PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid(7)                                                                        <= PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid(8)                                                                        <= PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid(9)                                                                        <= PriceSummaryWriter_l_inst_l_count_order_bus_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe(BUS_DATA_WIDTH/8 - 1 downto 0)                                           <= PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_strobe;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe(BUS_DATA_WIDTH/8 + BUS_DATA_WIDTH/8 - 1 downto BUS_DATA_WIDTH/8)         <= PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_strobe;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe(BUS_DATA_WIDTH/8 * 2 + BUS_DATA_WIDTH/8 - 1 downto BUS_DATA_WIDTH/8 * 2) <= PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_strobe;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe(BUS_DATA_WIDTH/8 * 3 + BUS_DATA_WIDTH/8 - 1 downto BUS_DATA_WIDTH/8 * 3) <= PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_strobe;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe(BUS_DATA_WIDTH/8 * 4 + BUS_DATA_WIDTH/8 - 1 downto BUS_DATA_WIDTH/8 * 4) <= PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_strobe;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe(BUS_DATA_WIDTH/8 * 5 + BUS_DATA_WIDTH/8 - 1 downto BUS_DATA_WIDTH/8 * 5) <= PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_strobe;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe(BUS_DATA_WIDTH/8 * 6 + BUS_DATA_WIDTH/8 - 1 downto BUS_DATA_WIDTH/8 * 6) <= PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_strobe;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe(BUS_DATA_WIDTH/8 * 7 + BUS_DATA_WIDTH/8 - 1 downto BUS_DATA_WIDTH/8 * 7) <= PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_strobe;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe(BUS_DATA_WIDTH/8 * 8 + BUS_DATA_WIDTH/8 - 1 downto BUS_DATA_WIDTH/8 * 8) <= PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_strobe;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe(BUS_DATA_WIDTH/8 * 9 + BUS_DATA_WIDTH/8 - 1 downto BUS_DATA_WIDTH/8 * 9) <= PriceSummaryWriter_l_inst_l_count_order_bus_wdat_strobe;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last(0)                                                                         <= PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_last;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last(1)                                                                         <= PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_last;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last(2)                                                                         <= PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_last;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last(3)                                                                         <= PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_last;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last(4)                                                                         <= PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_last;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last(5)                                                                         <= PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_last;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last(6)                                                                         <= PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_last;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last(7)                                                                         <= PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_last;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last(8)                                                                         <= PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_last;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last(9)                                                                         <= PriceSummaryWriter_l_inst_l_count_order_bus_wdat_last;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data(BUS_DATA_WIDTH - 1 downto 0)                                               <= PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_data;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data(BUS_DATA_WIDTH + BUS_DATA_WIDTH - 1 downto BUS_DATA_WIDTH)                 <= PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_data;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data(BUS_DATA_WIDTH * 2 + BUS_DATA_WIDTH - 1 downto BUS_DATA_WIDTH * 2)         <= PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_data;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data(BUS_DATA_WIDTH * 3 + BUS_DATA_WIDTH - 1 downto BUS_DATA_WIDTH * 3)         <= PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_data;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data(BUS_DATA_WIDTH * 4 + BUS_DATA_WIDTH - 1 downto BUS_DATA_WIDTH * 4)         <= PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_data;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data(BUS_DATA_WIDTH * 5 + BUS_DATA_WIDTH - 1 downto BUS_DATA_WIDTH * 5)         <= PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_data;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data(BUS_DATA_WIDTH * 6 + BUS_DATA_WIDTH - 1 downto BUS_DATA_WIDTH * 6)         <= PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_data;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data(BUS_DATA_WIDTH * 7 + BUS_DATA_WIDTH - 1 downto BUS_DATA_WIDTH * 7)         <= PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_data;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data(BUS_DATA_WIDTH * 8 + BUS_DATA_WIDTH - 1 downto BUS_DATA_WIDTH * 8)         <= PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_data;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data(BUS_DATA_WIDTH * 9 + BUS_DATA_WIDTH - 1 downto BUS_DATA_WIDTH * 9)         <= PriceSummaryWriter_l_inst_l_count_order_bus_wdat_data;
  PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_ready                                                                  <= WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready(2);
  PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_ready                                                                  <= WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready(2);
  PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_ready                                                           <= WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready(4);
  PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_ready                                                           <= WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready(4);
  PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_ready                                                               <= WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready(5);
  PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_ready                                                               <= WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready(5);
  PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_ready                                                           <= WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready(3);
  PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_ready                                                           <= WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready(3);
  PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_ready                                                             <= WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready(0);
  PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_ready                                                             <= WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready(0);
  PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_ready                                                             <= WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready(1);
  PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_ready                                                             <= WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready(1);
  PriceSummaryWriter_l_inst_l_count_order_bus_wreq_ready                                                              <= WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready(9);
  PriceSummaryWriter_l_inst_l_count_order_bus_wdat_ready                                                              <= WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready(9);
  PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_ready                                                                  <= WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready(6);
  PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_ready                                                                  <= WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready(6);
  PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_ready                                                                <= WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready(7);
  PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_ready                                                                <= WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready(7);
  PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_ready                                                                 <= WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready(8);
  PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_ready                                                                 <= WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready(8);
  RDAW64DW512LW8BS1BM16_inst : BusReadArbiterVec
  generic map(
    BUS_ADDR_WIDTH  => BUS_ADDR_WIDTH,
    BUS_DATA_WIDTH  => BUS_DATA_WIDTH,
    BUS_LEN_WIDTH   => BUS_LEN_WIDTH,
    NUM_SLAVE_PORTS => 7,
    ARB_METHOD      => "RR-STICKY",
    MAX_OUTSTANDING => 4,
    RAM_CONFIG      => "",
    SLV_REQ_SLICES  => true,
    MST_REQ_SLICE   => true,
    MST_DAT_SLICE   => true,
    SLV_DAT_SLICES  => true
  )
  port map(
    bcd_clk        => bcd_clk,
    bcd_reset      => bcd_reset,
    mst_rreq_valid => RDAW64DW512LW8BS1BM16_inst_mst_rreq_valid,
    mst_rreq_ready => RDAW64DW512LW8BS1BM16_inst_mst_rreq_ready,
    mst_rreq_addr  => RDAW64DW512LW8BS1BM16_inst_mst_rreq_addr,
    mst_rreq_len   => RDAW64DW512LW8BS1BM16_inst_mst_rreq_len,
    mst_rdat_valid => RDAW64DW512LW8BS1BM16_inst_mst_rdat_valid,
    mst_rdat_ready => RDAW64DW512LW8BS1BM16_inst_mst_rdat_ready,
    mst_rdat_data  => RDAW64DW512LW8BS1BM16_inst_mst_rdat_data,
    mst_rdat_last  => RDAW64DW512LW8BS1BM16_inst_mst_rdat_last,
    bsv_rreq_valid => RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid,
    bsv_rreq_ready => RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready,
    bsv_rreq_len   => RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len,
    bsv_rreq_addr  => RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr,
    bsv_rdat_valid => RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid,
    bsv_rdat_ready => RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready,
    bsv_rdat_last  => RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last,
    bsv_rdat_data  => RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data
  );

  rd_mst_rreq_valid                                                                                           <= RDAW64DW512LW8BS1BM16_inst_mst_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_mst_rreq_ready                                                                   <= rd_mst_rreq_ready;
  rd_mst_rreq_addr                                                                                            <= RDAW64DW512LW8BS1BM16_inst_mst_rreq_addr;
  rd_mst_rreq_len                                                                                             <= RDAW64DW512LW8BS1BM16_inst_mst_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_mst_rdat_valid                                                                   <= rd_mst_rdat_valid;
  rd_mst_rdat_ready                                                                                           <= RDAW64DW512LW8BS1BM16_inst_mst_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_mst_rdat_data                                                                    <= rd_mst_rdat_data;
  RDAW64DW512LW8BS1BM16_inst_mst_rdat_last                                                                    <= rd_mst_rdat_last;

  PriceSummary_Nucleus_inst_mmio_awvalid                                                                      <= mmio_awvalid;
  mmio_awready                                                                                                <= PriceSummary_Nucleus_inst_mmio_awready;
  PriceSummary_Nucleus_inst_mmio_awaddr                                                                       <= mmio_awaddr;
  PriceSummary_Nucleus_inst_mmio_wvalid                                                                       <= mmio_wvalid;
  mmio_wready                                                                                                 <= PriceSummary_Nucleus_inst_mmio_wready;
  PriceSummary_Nucleus_inst_mmio_wdata                                                                        <= mmio_wdata;
  PriceSummary_Nucleus_inst_mmio_wstrb                                                                        <= mmio_wstrb;
  mmio_bvalid                                                                                                 <= PriceSummary_Nucleus_inst_mmio_bvalid;
  PriceSummary_Nucleus_inst_mmio_bready                                                                       <= mmio_bready;
  mmio_bresp                                                                                                  <= PriceSummary_Nucleus_inst_mmio_bresp;
  PriceSummary_Nucleus_inst_mmio_arvalid                                                                      <= mmio_arvalid;
  mmio_arready                                                                                                <= PriceSummary_Nucleus_inst_mmio_arready;
  PriceSummary_Nucleus_inst_mmio_araddr                                                                       <= mmio_araddr;
  mmio_rvalid                                                                                                 <= PriceSummary_Nucleus_inst_mmio_rvalid;
  PriceSummary_Nucleus_inst_mmio_rready                                                                       <= mmio_rready;
  mmio_rdata                                                                                                  <= PriceSummary_Nucleus_inst_mmio_rdata;
  mmio_rresp                                                                                                  <= PriceSummary_Nucleus_inst_mmio_rresp;

  PriceSummary_Nucleus_inst_l_quantity_valid                                                                  <= PriceSummary_l_inst_l_quantity_valid;
  PriceSummary_l_inst_l_quantity_ready                                                                        <= PriceSummary_Nucleus_inst_l_quantity_ready;
  PriceSummary_Nucleus_inst_l_quantity_dvalid                                                                 <= PriceSummary_l_inst_l_quantity_dvalid;
  PriceSummary_Nucleus_inst_l_quantity_last                                                                   <= PriceSummary_l_inst_l_quantity_last;
  PriceSummary_Nucleus_inst_l_quantity                                                                        <= PriceSummary_l_inst_l_quantity;

  PriceSummary_Nucleus_inst_l_extendedprice_valid                                                             <= PriceSummary_l_inst_l_extendedprice_valid;
  PriceSummary_l_inst_l_extendedprice_ready                                                                   <= PriceSummary_Nucleus_inst_l_extendedprice_ready;
  PriceSummary_Nucleus_inst_l_extendedprice_dvalid                                                            <= PriceSummary_l_inst_l_extendedprice_dvalid;
  PriceSummary_Nucleus_inst_l_extendedprice_last                                                              <= PriceSummary_l_inst_l_extendedprice_last;
  PriceSummary_Nucleus_inst_l_extendedprice                                                                   <= PriceSummary_l_inst_l_extendedprice;

  PriceSummary_Nucleus_inst_l_discount_valid                                                                  <= PriceSummary_l_inst_l_discount_valid;
  PriceSummary_l_inst_l_discount_ready                                                                        <= PriceSummary_Nucleus_inst_l_discount_ready;
  PriceSummary_Nucleus_inst_l_discount_dvalid                                                                 <= PriceSummary_l_inst_l_discount_dvalid;
  PriceSummary_Nucleus_inst_l_discount_last                                                                   <= PriceSummary_l_inst_l_discount_last;
  PriceSummary_Nucleus_inst_l_discount                                                                        <= PriceSummary_l_inst_l_discount;

  PriceSummary_Nucleus_inst_l_tax_valid                                                                       <= PriceSummary_l_inst_l_tax_valid;
  PriceSummary_l_inst_l_tax_ready                                                                             <= PriceSummary_Nucleus_inst_l_tax_ready;
  PriceSummary_Nucleus_inst_l_tax_dvalid                                                                      <= PriceSummary_l_inst_l_tax_dvalid;
  PriceSummary_Nucleus_inst_l_tax_last                                                                        <= PriceSummary_l_inst_l_tax_last;
  PriceSummary_Nucleus_inst_l_tax                                                                             <= PriceSummary_l_inst_l_tax;

  PriceSummary_Nucleus_inst_l_returnflag_valid                                                                <= PriceSummary_l_inst_l_returnflag_valid;
  PriceSummary_l_inst_l_returnflag_ready                                                                      <= PriceSummary_Nucleus_inst_l_returnflag_ready;
  PriceSummary_Nucleus_inst_l_returnflag_dvalid                                                               <= PriceSummary_l_inst_l_returnflag_dvalid;
  PriceSummary_Nucleus_inst_l_returnflag_last                                                                 <= PriceSummary_l_inst_l_returnflag_last;
  PriceSummary_Nucleus_inst_l_returnflag_length                                                               <= PriceSummary_l_inst_l_returnflag_length;
  PriceSummary_Nucleus_inst_l_returnflag_count                                                                <= PriceSummary_l_inst_l_returnflag_count;
  PriceSummary_Nucleus_inst_l_returnflag_chars_valid                                                          <= PriceSummary_l_inst_l_returnflag_chars_valid;
  PriceSummary_l_inst_l_returnflag_chars_ready                                                                <= PriceSummary_Nucleus_inst_l_returnflag_chars_ready;
  PriceSummary_Nucleus_inst_l_returnflag_chars_dvalid                                                         <= PriceSummary_l_inst_l_returnflag_chars_dvalid;
  PriceSummary_Nucleus_inst_l_returnflag_chars_last                                                           <= PriceSummary_l_inst_l_returnflag_chars_last;
  PriceSummary_Nucleus_inst_l_returnflag_chars                                                                <= PriceSummary_l_inst_l_returnflag_chars;
  PriceSummary_Nucleus_inst_l_returnflag_chars_count                                                          <= PriceSummary_l_inst_l_returnflag_chars_count;

  PriceSummary_Nucleus_inst_l_linestatus_valid                                                                <= PriceSummary_l_inst_l_linestatus_valid;
  PriceSummary_l_inst_l_linestatus_ready                                                                      <= PriceSummary_Nucleus_inst_l_linestatus_ready;
  PriceSummary_Nucleus_inst_l_linestatus_dvalid                                                               <= PriceSummary_l_inst_l_linestatus_dvalid;
  PriceSummary_Nucleus_inst_l_linestatus_last                                                                 <= PriceSummary_l_inst_l_linestatus_last;
  PriceSummary_Nucleus_inst_l_linestatus_length                                                               <= PriceSummary_l_inst_l_linestatus_length;
  PriceSummary_Nucleus_inst_l_linestatus_count                                                                <= PriceSummary_l_inst_l_linestatus_count;
  PriceSummary_Nucleus_inst_l_linestatus_chars_valid                                                          <= PriceSummary_l_inst_l_linestatus_chars_valid;
  PriceSummary_l_inst_l_linestatus_chars_ready                                                                <= PriceSummary_Nucleus_inst_l_linestatus_chars_ready;
  PriceSummary_Nucleus_inst_l_linestatus_chars_dvalid                                                         <= PriceSummary_l_inst_l_linestatus_chars_dvalid;
  PriceSummary_Nucleus_inst_l_linestatus_chars_last                                                           <= PriceSummary_l_inst_l_linestatus_chars_last;
  PriceSummary_Nucleus_inst_l_linestatus_chars                                                                <= PriceSummary_l_inst_l_linestatus_chars;
  PriceSummary_Nucleus_inst_l_linestatus_chars_count                                                          <= PriceSummary_l_inst_l_linestatus_chars_count;

  PriceSummary_Nucleus_inst_l_shipdate_valid                                                                  <= PriceSummary_l_inst_l_shipdate_valid;
  PriceSummary_l_inst_l_shipdate_ready                                                                        <= PriceSummary_Nucleus_inst_l_shipdate_ready;
  PriceSummary_Nucleus_inst_l_shipdate_dvalid                                                                 <= PriceSummary_l_inst_l_shipdate_dvalid;
  PriceSummary_Nucleus_inst_l_shipdate_last                                                                   <= PriceSummary_l_inst_l_shipdate_last;
  PriceSummary_Nucleus_inst_l_shipdate                                                                        <= PriceSummary_l_inst_l_shipdate;

  PriceSummary_Nucleus_inst_l_quantity_unl_valid                                                              <= PriceSummary_l_inst_l_quantity_unl_valid;
  PriceSummary_l_inst_l_quantity_unl_ready                                                                    <= PriceSummary_Nucleus_inst_l_quantity_unl_ready;
  PriceSummary_Nucleus_inst_l_quantity_unl_tag                                                                <= PriceSummary_l_inst_l_quantity_unl_tag;

  PriceSummary_Nucleus_inst_l_extendedprice_unl_valid                                                         <= PriceSummary_l_inst_l_extendedprice_unl_valid;
  PriceSummary_l_inst_l_extendedprice_unl_ready                                                               <= PriceSummary_Nucleus_inst_l_extendedprice_unl_ready;
  PriceSummary_Nucleus_inst_l_extendedprice_unl_tag                                                           <= PriceSummary_l_inst_l_extendedprice_unl_tag;

  PriceSummary_Nucleus_inst_l_discount_unl_valid                                                              <= PriceSummary_l_inst_l_discount_unl_valid;
  PriceSummary_l_inst_l_discount_unl_ready                                                                    <= PriceSummary_Nucleus_inst_l_discount_unl_ready;
  PriceSummary_Nucleus_inst_l_discount_unl_tag                                                                <= PriceSummary_l_inst_l_discount_unl_tag;

  PriceSummary_Nucleus_inst_l_tax_unl_valid                                                                   <= PriceSummary_l_inst_l_tax_unl_valid;
  PriceSummary_l_inst_l_tax_unl_ready                                                                         <= PriceSummary_Nucleus_inst_l_tax_unl_ready;
  PriceSummary_Nucleus_inst_l_tax_unl_tag                                                                     <= PriceSummary_l_inst_l_tax_unl_tag;

  PriceSummary_Nucleus_inst_l_returnflag_unl_valid                                                            <= PriceSummary_l_inst_l_returnflag_unl_valid;
  PriceSummary_l_inst_l_returnflag_unl_ready                                                                  <= PriceSummary_Nucleus_inst_l_returnflag_unl_ready;
  PriceSummary_Nucleus_inst_l_returnflag_unl_tag                                                              <= PriceSummary_l_inst_l_returnflag_unl_tag;

  PriceSummary_Nucleus_inst_l_linestatus_unl_valid                                                            <= PriceSummary_l_inst_l_linestatus_unl_valid;
  PriceSummary_l_inst_l_linestatus_unl_ready                                                                  <= PriceSummary_Nucleus_inst_l_linestatus_unl_ready;
  PriceSummary_Nucleus_inst_l_linestatus_unl_tag                                                              <= PriceSummary_l_inst_l_linestatus_unl_tag;

  PriceSummary_Nucleus_inst_l_shipdate_unl_valid                                                              <= PriceSummary_l_inst_l_shipdate_unl_valid;
  PriceSummary_l_inst_l_shipdate_unl_ready                                                                    <= PriceSummary_Nucleus_inst_l_shipdate_unl_ready;
  PriceSummary_Nucleus_inst_l_shipdate_unl_tag                                                                <= PriceSummary_l_inst_l_shipdate_unl_tag;

  PriceSummary_l_inst_l_quantity_cmd_valid                                                                    <= PriceSummary_Nucleus_inst_l_quantity_cmd_valid;
  PriceSummary_Nucleus_inst_l_quantity_cmd_ready                                                              <= PriceSummary_l_inst_l_quantity_cmd_ready;
  PriceSummary_l_inst_l_quantity_cmd_firstIdx                                                                 <= PriceSummary_Nucleus_inst_l_quantity_cmd_firstIdx;
  PriceSummary_l_inst_l_quantity_cmd_lastIdx                                                                  <= PriceSummary_Nucleus_inst_l_quantity_cmd_lastIdx;
  PriceSummary_l_inst_l_quantity_cmd_ctrl                                                                     <= PriceSummary_Nucleus_inst_l_quantity_cmd_ctrl;
  PriceSummary_l_inst_l_quantity_cmd_tag                                                                      <= PriceSummary_Nucleus_inst_l_quantity_cmd_tag;

  PriceSummary_l_inst_l_extendedprice_cmd_valid                                                               <= PriceSummary_Nucleus_inst_l_extendedprice_cmd_valid;
  PriceSummary_Nucleus_inst_l_extendedprice_cmd_ready                                                         <= PriceSummary_l_inst_l_extendedprice_cmd_ready;
  PriceSummary_l_inst_l_extendedprice_cmd_firstIdx                                                            <= PriceSummary_Nucleus_inst_l_extendedprice_cmd_firstIdx;
  PriceSummary_l_inst_l_extendedprice_cmd_lastIdx                                                             <= PriceSummary_Nucleus_inst_l_extendedprice_cmd_lastIdx;
  PriceSummary_l_inst_l_extendedprice_cmd_ctrl                                                                <= PriceSummary_Nucleus_inst_l_extendedprice_cmd_ctrl;
  PriceSummary_l_inst_l_extendedprice_cmd_tag                                                                 <= PriceSummary_Nucleus_inst_l_extendedprice_cmd_tag;

  PriceSummary_l_inst_l_discount_cmd_valid                                                                    <= PriceSummary_Nucleus_inst_l_discount_cmd_valid;
  PriceSummary_Nucleus_inst_l_discount_cmd_ready                                                              <= PriceSummary_l_inst_l_discount_cmd_ready;
  PriceSummary_l_inst_l_discount_cmd_firstIdx                                                                 <= PriceSummary_Nucleus_inst_l_discount_cmd_firstIdx;
  PriceSummary_l_inst_l_discount_cmd_lastIdx                                                                  <= PriceSummary_Nucleus_inst_l_discount_cmd_lastIdx;
  PriceSummary_l_inst_l_discount_cmd_ctrl                                                                     <= PriceSummary_Nucleus_inst_l_discount_cmd_ctrl;
  PriceSummary_l_inst_l_discount_cmd_tag                                                                      <= PriceSummary_Nucleus_inst_l_discount_cmd_tag;

  PriceSummary_l_inst_l_tax_cmd_valid                                                                         <= PriceSummary_Nucleus_inst_l_tax_cmd_valid;
  PriceSummary_Nucleus_inst_l_tax_cmd_ready                                                                   <= PriceSummary_l_inst_l_tax_cmd_ready;
  PriceSummary_l_inst_l_tax_cmd_firstIdx                                                                      <= PriceSummary_Nucleus_inst_l_tax_cmd_firstIdx;
  PriceSummary_l_inst_l_tax_cmd_lastIdx                                                                       <= PriceSummary_Nucleus_inst_l_tax_cmd_lastIdx;
  PriceSummary_l_inst_l_tax_cmd_ctrl                                                                          <= PriceSummary_Nucleus_inst_l_tax_cmd_ctrl;
  PriceSummary_l_inst_l_tax_cmd_tag                                                                           <= PriceSummary_Nucleus_inst_l_tax_cmd_tag;

  PriceSummary_l_inst_l_returnflag_cmd_valid                                                                  <= PriceSummary_Nucleus_inst_l_returnflag_cmd_valid;
  PriceSummary_Nucleus_inst_l_returnflag_cmd_ready                                                            <= PriceSummary_l_inst_l_returnflag_cmd_ready;
  PriceSummary_l_inst_l_returnflag_cmd_firstIdx                                                               <= PriceSummary_Nucleus_inst_l_returnflag_cmd_firstIdx;
  PriceSummary_l_inst_l_returnflag_cmd_lastIdx                                                                <= PriceSummary_Nucleus_inst_l_returnflag_cmd_lastIdx;
  PriceSummary_l_inst_l_returnflag_cmd_ctrl                                                                   <= PriceSummary_Nucleus_inst_l_returnflag_cmd_ctrl;
  PriceSummary_l_inst_l_returnflag_cmd_tag                                                                    <= PriceSummary_Nucleus_inst_l_returnflag_cmd_tag;

  PriceSummary_l_inst_l_linestatus_cmd_valid                                                                  <= PriceSummary_Nucleus_inst_l_linestatus_cmd_valid;
  PriceSummary_Nucleus_inst_l_linestatus_cmd_ready                                                            <= PriceSummary_l_inst_l_linestatus_cmd_ready;
  PriceSummary_l_inst_l_linestatus_cmd_firstIdx                                                               <= PriceSummary_Nucleus_inst_l_linestatus_cmd_firstIdx;
  PriceSummary_l_inst_l_linestatus_cmd_lastIdx                                                                <= PriceSummary_Nucleus_inst_l_linestatus_cmd_lastIdx;
  PriceSummary_l_inst_l_linestatus_cmd_ctrl                                                                   <= PriceSummary_Nucleus_inst_l_linestatus_cmd_ctrl;
  PriceSummary_l_inst_l_linestatus_cmd_tag                                                                    <= PriceSummary_Nucleus_inst_l_linestatus_cmd_tag;

  PriceSummary_l_inst_l_shipdate_cmd_valid                                                                    <= PriceSummary_Nucleus_inst_l_shipdate_cmd_valid;
  PriceSummary_Nucleus_inst_l_shipdate_cmd_ready                                                              <= PriceSummary_l_inst_l_shipdate_cmd_ready;
  PriceSummary_l_inst_l_shipdate_cmd_firstIdx                                                                 <= PriceSummary_Nucleus_inst_l_shipdate_cmd_firstIdx;
  PriceSummary_l_inst_l_shipdate_cmd_lastIdx                                                                  <= PriceSummary_Nucleus_inst_l_shipdate_cmd_lastIdx;
  PriceSummary_l_inst_l_shipdate_cmd_ctrl                                                                     <= PriceSummary_Nucleus_inst_l_shipdate_cmd_ctrl;
  PriceSummary_l_inst_l_shipdate_cmd_tag                                                                      <= PriceSummary_Nucleus_inst_l_shipdate_cmd_tag;

  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(0)                                                                <= PriceSummary_l_inst_l_quantity_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(1)                                                                <= PriceSummary_l_inst_l_extendedprice_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(2)                                                                <= PriceSummary_l_inst_l_discount_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(3)                                                                <= PriceSummary_l_inst_l_tax_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(4)                                                                <= PriceSummary_l_inst_l_returnflag_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(5)                                                                <= PriceSummary_l_inst_l_linestatus_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(6)                                                                <= PriceSummary_l_inst_l_shipdate_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH - 1 downto 0)                                         <= PriceSummary_l_inst_l_quantity_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH + BUS_LEN_WIDTH - 1 downto BUS_LEN_WIDTH)             <= PriceSummary_l_inst_l_extendedprice_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH * 2 + BUS_LEN_WIDTH - 1 downto BUS_LEN_WIDTH * 2)     <= PriceSummary_l_inst_l_discount_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH * 3 + BUS_LEN_WIDTH - 1 downto BUS_LEN_WIDTH * 3)     <= PriceSummary_l_inst_l_tax_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH * 4 + BUS_LEN_WIDTH - 1 downto BUS_LEN_WIDTH * 4)     <= PriceSummary_l_inst_l_returnflag_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH * 5 + BUS_LEN_WIDTH - 1 downto BUS_LEN_WIDTH * 5)     <= PriceSummary_l_inst_l_linestatus_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH * 6 + BUS_LEN_WIDTH - 1 downto BUS_LEN_WIDTH * 6)     <= PriceSummary_l_inst_l_shipdate_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH - 1 downto 0)                                       <= PriceSummary_l_inst_l_quantity_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH + BUS_ADDR_WIDTH - 1 downto BUS_ADDR_WIDTH)         <= PriceSummary_l_inst_l_extendedprice_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH * 2 + BUS_ADDR_WIDTH - 1 downto BUS_ADDR_WIDTH * 2) <= PriceSummary_l_inst_l_discount_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH * 3 + BUS_ADDR_WIDTH - 1 downto BUS_ADDR_WIDTH * 3) <= PriceSummary_l_inst_l_tax_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH * 4 + BUS_ADDR_WIDTH - 1 downto BUS_ADDR_WIDTH * 4) <= PriceSummary_l_inst_l_returnflag_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH * 5 + BUS_ADDR_WIDTH - 1 downto BUS_ADDR_WIDTH * 5) <= PriceSummary_l_inst_l_linestatus_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH * 6 + BUS_ADDR_WIDTH - 1 downto BUS_ADDR_WIDTH * 6) <= PriceSummary_l_inst_l_shipdate_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(0)                                                                <= PriceSummary_l_inst_l_quantity_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(1)                                                                <= PriceSummary_l_inst_l_extendedprice_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(2)                                                                <= PriceSummary_l_inst_l_discount_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(3)                                                                <= PriceSummary_l_inst_l_tax_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(4)                                                                <= PriceSummary_l_inst_l_returnflag_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(5)                                                                <= PriceSummary_l_inst_l_linestatus_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(6)                                                                <= PriceSummary_l_inst_l_shipdate_bus_rdat_ready;
  PriceSummary_l_inst_l_tax_bus_rreq_ready                                                                    <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(3);
  PriceSummary_l_inst_l_tax_bus_rdat_valid                                                                    <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(3);
  PriceSummary_l_inst_l_tax_bus_rdat_last                                                                     <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(3);
  PriceSummary_l_inst_l_tax_bus_rdat_data                                                                     <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH * 3 + BUS_DATA_WIDTH - 1 downto BUS_DATA_WIDTH * 3);
  PriceSummary_l_inst_l_shipdate_bus_rreq_ready                                                               <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(6);
  PriceSummary_l_inst_l_shipdate_bus_rdat_valid                                                               <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(6);
  PriceSummary_l_inst_l_shipdate_bus_rdat_last                                                                <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(6);
  PriceSummary_l_inst_l_shipdate_bus_rdat_data                                                                <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH * 6 + BUS_DATA_WIDTH - 1 downto BUS_DATA_WIDTH * 6);
  PriceSummary_l_inst_l_returnflag_bus_rreq_ready                                                             <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(4);
  PriceSummary_l_inst_l_returnflag_bus_rdat_valid                                                             <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(4);
  PriceSummary_l_inst_l_returnflag_bus_rdat_last                                                              <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(4);
  PriceSummary_l_inst_l_returnflag_bus_rdat_data                                                              <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH * 4 + BUS_DATA_WIDTH - 1 downto BUS_DATA_WIDTH * 4);
  PriceSummary_l_inst_l_quantity_bus_rreq_ready                                                               <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(0);
  PriceSummary_l_inst_l_quantity_bus_rdat_valid                                                               <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(0);
  PriceSummary_l_inst_l_quantity_bus_rdat_last                                                                <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(0);
  PriceSummary_l_inst_l_quantity_bus_rdat_data                                                                <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH - 1 downto 0);
  PriceSummary_l_inst_l_linestatus_bus_rreq_ready                                                             <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(5);
  PriceSummary_l_inst_l_linestatus_bus_rdat_valid                                                             <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(5);
  PriceSummary_l_inst_l_linestatus_bus_rdat_last                                                              <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(5);
  PriceSummary_l_inst_l_linestatus_bus_rdat_data                                                              <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH * 5 + BUS_DATA_WIDTH - 1 downto BUS_DATA_WIDTH * 5);
  PriceSummary_l_inst_l_extendedprice_bus_rreq_ready                                                          <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(1);
  PriceSummary_l_inst_l_extendedprice_bus_rdat_valid                                                          <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(1);
  PriceSummary_l_inst_l_extendedprice_bus_rdat_last                                                           <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(1);
  PriceSummary_l_inst_l_extendedprice_bus_rdat_data                                                           <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH + BUS_DATA_WIDTH - 1 downto BUS_DATA_WIDTH);
  PriceSummary_l_inst_l_discount_bus_rreq_ready                                                               <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(2);
  PriceSummary_l_inst_l_discount_bus_rdat_valid                                                               <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(2);
  PriceSummary_l_inst_l_discount_bus_rdat_last                                                                <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(2);
  PriceSummary_l_inst_l_discount_bus_rdat_data                                                                <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH * 2 + BUS_DATA_WIDTH - 1 downto BUS_DATA_WIDTH * 2);

end architecture;