-- Copyright 2018-2019 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
-- This file was generated by Fletchgen. Modify this file at your own risk.

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

LIBRARY work;
USE work.Array_pkg.ALL;
USE work.mmio_pkg.ALL;

ENTITY PriceSummary_Nucleus IS
  GENERIC (
    INDEX_WIDTH : INTEGER := 32;
    TAG_WIDTH : INTEGER := 1;
    L_QUANTITY_BUS_ADDR_WIDTH : INTEGER := 64;
    L_EXTENDEDPRICE_BUS_ADDR_WIDTH : INTEGER := 64;
    L_DISCOUNT_BUS_ADDR_WIDTH : INTEGER := 64;
    L_TAX_BUS_ADDR_WIDTH : INTEGER := 64;
    L_RETURNFLAG_BUS_ADDR_WIDTH : INTEGER := 64;
    L_LINESTATUS_BUS_ADDR_WIDTH : INTEGER := 64;
    L_SHIPDATE_BUS_ADDR_WIDTH : INTEGER := 64;
    L_RETURNFLAG_O_BUS_ADDR_WIDTH : INTEGER := 64;
    L_LINESTATUS_O_BUS_ADDR_WIDTH : INTEGER := 64;
    L_SUM_QTY_BUS_ADDR_WIDTH : INTEGER := 64;
    L_SUM_BASE_PRICE_BUS_ADDR_WIDTH : INTEGER := 64;
    L_SUM_DISC_PRICE_BUS_ADDR_WIDTH : INTEGER := 64;
    L_SUM_CHARGE_BUS_ADDR_WIDTH : INTEGER := 64;
    L_AVG_QTY_BUS_ADDR_WIDTH : INTEGER := 64;
    L_AVG_PRICE_BUS_ADDR_WIDTH : INTEGER := 64;
    L_AVG_DISC_BUS_ADDR_WIDTH : INTEGER := 64;
    L_COUNT_ORDER_BUS_ADDR_WIDTH : INTEGER := 64
  );
  PORT (
    kcd_clk : IN STD_LOGIC;
    kcd_reset : IN STD_LOGIC;
    mmio_awvalid : IN STD_LOGIC;
    mmio_awready : OUT STD_LOGIC;
    mmio_awaddr : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    mmio_wvalid : IN STD_LOGIC;
    mmio_wready : OUT STD_LOGIC;
    mmio_wdata : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    mmio_wstrb : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    mmio_bvalid : OUT STD_LOGIC;
    mmio_bready : IN STD_LOGIC;
    mmio_bresp : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    mmio_arvalid : IN STD_LOGIC;
    mmio_arready : OUT STD_LOGIC;
    mmio_araddr : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    mmio_rvalid : OUT STD_LOGIC;
    mmio_rready : IN STD_LOGIC;
    mmio_rdata : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    mmio_rresp : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    l_quantity_valid : IN STD_LOGIC;
    l_quantity_ready : OUT STD_LOGIC;
    l_quantity_dvalid : IN STD_LOGIC;
    l_quantity_last : IN STD_LOGIC;
    l_quantity : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
    l_extendedprice_valid : IN STD_LOGIC;
    l_extendedprice_ready : OUT STD_LOGIC;
    l_extendedprice_dvalid : IN STD_LOGIC;
    l_extendedprice_last : IN STD_LOGIC;
    l_extendedprice : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
    l_discount_valid : IN STD_LOGIC;
    l_discount_ready : OUT STD_LOGIC;
    l_discount_dvalid : IN STD_LOGIC;
    l_discount_last : IN STD_LOGIC;
    l_discount : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
    l_tax_valid : IN STD_LOGIC;
    l_tax_ready : OUT STD_LOGIC;
    l_tax_dvalid : IN STD_LOGIC;
    l_tax_last : IN STD_LOGIC;
    l_tax : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
    l_returnflag_valid : IN STD_LOGIC;
    l_returnflag_ready : OUT STD_LOGIC;
    l_returnflag_dvalid : IN STD_LOGIC;
    l_returnflag_last : IN STD_LOGIC;
    l_returnflag_length : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    l_returnflag_count : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    l_returnflag_chars_valid : IN STD_LOGIC;
    l_returnflag_chars_ready : OUT STD_LOGIC;
    l_returnflag_chars_dvalid : IN STD_LOGIC;
    l_returnflag_chars_last : IN STD_LOGIC;
    l_returnflag_chars : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    l_returnflag_chars_count : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    l_linestatus_valid : IN STD_LOGIC;
    l_linestatus_ready : OUT STD_LOGIC;
    l_linestatus_dvalid : IN STD_LOGIC;
    l_linestatus_last : IN STD_LOGIC;
    l_linestatus_length : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    l_linestatus_count : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    l_linestatus_chars_valid : IN STD_LOGIC;
    l_linestatus_chars_ready : OUT STD_LOGIC;
    l_linestatus_chars_dvalid : IN STD_LOGIC;
    l_linestatus_chars_last : IN STD_LOGIC;
    l_linestatus_chars : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
    l_linestatus_chars_count : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
    l_shipdate_valid : IN STD_LOGIC;
    l_shipdate_ready : OUT STD_LOGIC;
    l_shipdate_dvalid : IN STD_LOGIC;
    l_shipdate_last : IN STD_LOGIC;
    l_shipdate : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    l_quantity_unl_valid : IN STD_LOGIC;
    l_quantity_unl_ready : OUT STD_LOGIC;
    l_quantity_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
    l_extendedprice_unl_valid : IN STD_LOGIC;
    l_extendedprice_unl_ready : OUT STD_LOGIC;
    l_extendedprice_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
    l_discount_unl_valid : IN STD_LOGIC;
    l_discount_unl_ready : OUT STD_LOGIC;
    l_discount_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
    l_tax_unl_valid : IN STD_LOGIC;
    l_tax_unl_ready : OUT STD_LOGIC;
    l_tax_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
    l_returnflag_unl_valid : IN STD_LOGIC;
    l_returnflag_unl_ready : OUT STD_LOGIC;
    l_returnflag_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
    l_linestatus_unl_valid : IN STD_LOGIC;
    l_linestatus_unl_ready : OUT STD_LOGIC;
    l_linestatus_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
    l_shipdate_unl_valid : IN STD_LOGIC;
    l_shipdate_unl_ready : OUT STD_LOGIC;
    l_shipdate_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
    l_quantity_cmd_valid : OUT STD_LOGIC;
    l_quantity_cmd_ready : IN STD_LOGIC;
    l_quantity_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
    l_quantity_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
    l_quantity_cmd_ctrl : OUT STD_LOGIC_VECTOR(L_QUANTITY_BUS_ADDR_WIDTH - 1 DOWNTO 0);
    l_quantity_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
    l_extendedprice_cmd_valid : OUT STD_LOGIC;
    l_extendedprice_cmd_ready : IN STD_LOGIC;
    l_extendedprice_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
    l_extendedprice_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
    l_extendedprice_cmd_ctrl : OUT STD_LOGIC_VECTOR(L_EXTENDEDPRICE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
    l_extendedprice_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
    l_discount_cmd_valid : OUT STD_LOGIC;
    l_discount_cmd_ready : IN STD_LOGIC;
    l_discount_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
    l_discount_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
    l_discount_cmd_ctrl : OUT STD_LOGIC_VECTOR(L_DISCOUNT_BUS_ADDR_WIDTH - 1 DOWNTO 0);
    l_discount_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
    l_tax_cmd_valid : OUT STD_LOGIC;
    l_tax_cmd_ready : IN STD_LOGIC;
    l_tax_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
    l_tax_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
    l_tax_cmd_ctrl : OUT STD_LOGIC_VECTOR(L_TAX_BUS_ADDR_WIDTH - 1 DOWNTO 0);
    l_tax_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
    l_returnflag_cmd_valid : OUT STD_LOGIC;
    l_returnflag_cmd_ready : IN STD_LOGIC;
    l_returnflag_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
    l_returnflag_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
    l_returnflag_cmd_ctrl : OUT STD_LOGIC_VECTOR(L_RETURNFLAG_BUS_ADDR_WIDTH * 2 - 1 DOWNTO 0);
    l_returnflag_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
    l_linestatus_cmd_valid : OUT STD_LOGIC;
    l_linestatus_cmd_ready : IN STD_LOGIC;
    l_linestatus_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
    l_linestatus_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
    l_linestatus_cmd_ctrl : OUT STD_LOGIC_VECTOR(L_LINESTATUS_BUS_ADDR_WIDTH * 2 - 1 DOWNTO 0);
    l_linestatus_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
    l_shipdate_cmd_valid : OUT STD_LOGIC;
    l_shipdate_cmd_ready : IN STD_LOGIC;
    l_shipdate_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
    l_shipdate_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
    l_shipdate_cmd_ctrl : OUT STD_LOGIC_VECTOR(L_SHIPDATE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
    l_shipdate_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
    l_returnflag_o_valid : OUT STD_LOGIC;
    l_returnflag_o_ready : IN STD_LOGIC;
    l_returnflag_o_dvalid : OUT STD_LOGIC;
    l_returnflag_o_last : OUT STD_LOGIC;
    l_returnflag_o_length : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    l_returnflag_o_count : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
    l_returnflag_o_chars_valid : OUT STD_LOGIC;
    l_returnflag_o_chars_ready : IN STD_LOGIC;
    l_returnflag_o_chars_dvalid : OUT STD_LOGIC;
    l_returnflag_o_chars_last : OUT STD_LOGIC;
    l_returnflag_o_chars : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    l_returnflag_o_chars_count : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
    l_linestatus_o_valid : OUT STD_LOGIC;
    l_linestatus_o_ready : IN STD_LOGIC;
    l_linestatus_o_dvalid : OUT STD_LOGIC;
    l_linestatus_o_last : OUT STD_LOGIC;
    l_linestatus_o_length : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    l_linestatus_o_count : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
    l_linestatus_o_chars_valid : OUT STD_LOGIC;
    l_linestatus_o_chars_ready : IN STD_LOGIC;
    l_linestatus_o_chars_dvalid : OUT STD_LOGIC;
    l_linestatus_o_chars_last : OUT STD_LOGIC;
    l_linestatus_o_chars : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
    l_linestatus_o_chars_count : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
    l_sum_qty_valid : OUT STD_LOGIC;
    l_sum_qty_ready : IN STD_LOGIC;
    l_sum_qty_dvalid : OUT STD_LOGIC;
    l_sum_qty_last : OUT STD_LOGIC;
    l_sum_qty : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
    l_sum_base_price_valid : OUT STD_LOGIC;
    l_sum_base_price_ready : IN STD_LOGIC;
    l_sum_base_price_dvalid : OUT STD_LOGIC;
    l_sum_base_price_last : OUT STD_LOGIC;
    l_sum_base_price : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
    l_sum_disc_price_valid : OUT STD_LOGIC;
    l_sum_disc_price_ready : IN STD_LOGIC;
    l_sum_disc_price_dvalid : OUT STD_LOGIC;
    l_sum_disc_price_last : OUT STD_LOGIC;
    l_sum_disc_price : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
    l_sum_charge_valid : OUT STD_LOGIC;
    l_sum_charge_ready : IN STD_LOGIC;
    l_sum_charge_dvalid : OUT STD_LOGIC;
    l_sum_charge_last : OUT STD_LOGIC;
    l_sum_charge : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
    l_avg_qty_valid : OUT STD_LOGIC;
    l_avg_qty_ready : IN STD_LOGIC;
    l_avg_qty_dvalid : OUT STD_LOGIC;
    l_avg_qty_last : OUT STD_LOGIC;
    l_avg_qty : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
    l_avg_price_valid : OUT STD_LOGIC;
    l_avg_price_ready : IN STD_LOGIC;
    l_avg_price_dvalid : OUT STD_LOGIC;
    l_avg_price_last : OUT STD_LOGIC;
    l_avg_price : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
    l_avg_disc_valid : OUT STD_LOGIC;
    l_avg_disc_ready : IN STD_LOGIC;
    l_avg_disc_dvalid : OUT STD_LOGIC;
    l_avg_disc_last : OUT STD_LOGIC;
    l_avg_disc : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
    l_count_order_valid : OUT STD_LOGIC;
    l_count_order_ready : IN STD_LOGIC;
    l_count_order_dvalid : OUT STD_LOGIC;
    l_count_order_last : OUT STD_LOGIC;
    l_count_order : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
    l_returnflag_o_unl_valid : IN STD_LOGIC;
    l_returnflag_o_unl_ready : OUT STD_LOGIC;
    l_returnflag_o_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
    l_linestatus_o_unl_valid : IN STD_LOGIC;
    l_linestatus_o_unl_ready : OUT STD_LOGIC;
    l_linestatus_o_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
    l_sum_qty_unl_valid : IN STD_LOGIC;
    l_sum_qty_unl_ready : OUT STD_LOGIC;
    l_sum_qty_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
    l_sum_base_price_unl_valid : IN STD_LOGIC;
    l_sum_base_price_unl_ready : OUT STD_LOGIC;
    l_sum_base_price_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
    l_sum_disc_price_unl_valid : IN STD_LOGIC;
    l_sum_disc_price_unl_ready : OUT STD_LOGIC;
    l_sum_disc_price_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
    l_sum_charge_unl_valid : IN STD_LOGIC;
    l_sum_charge_unl_ready : OUT STD_LOGIC;
    l_sum_charge_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
    l_avg_qty_unl_valid : IN STD_LOGIC;
    l_avg_qty_unl_ready : OUT STD_LOGIC;
    l_avg_qty_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
    l_avg_price_unl_valid : IN STD_LOGIC;
    l_avg_price_unl_ready : OUT STD_LOGIC;
    l_avg_price_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
    l_avg_disc_unl_valid : IN STD_LOGIC;
    l_avg_disc_unl_ready : OUT STD_LOGIC;
    l_avg_disc_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
    l_count_order_unl_valid : IN STD_LOGIC;
    l_count_order_unl_ready : OUT STD_LOGIC;
    l_count_order_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
    l_returnflag_o_cmd_valid : OUT STD_LOGIC;
    l_returnflag_o_cmd_ready : IN STD_LOGIC;
    l_returnflag_o_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
    l_returnflag_o_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
    l_returnflag_o_cmd_ctrl : OUT STD_LOGIC_VECTOR(L_RETURNFLAG_O_BUS_ADDR_WIDTH * 2 - 1 DOWNTO 0);
    l_returnflag_o_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
    l_linestatus_o_cmd_valid : OUT STD_LOGIC;
    l_linestatus_o_cmd_ready : IN STD_LOGIC;
    l_linestatus_o_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
    l_linestatus_o_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
    l_linestatus_o_cmd_ctrl : OUT STD_LOGIC_VECTOR(L_LINESTATUS_O_BUS_ADDR_WIDTH * 2 - 1 DOWNTO 0);
    l_linestatus_o_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
    l_sum_qty_cmd_valid : OUT STD_LOGIC;
    l_sum_qty_cmd_ready : IN STD_LOGIC;
    l_sum_qty_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
    l_sum_qty_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
    l_sum_qty_cmd_ctrl : OUT STD_LOGIC_VECTOR(L_SUM_QTY_BUS_ADDR_WIDTH - 1 DOWNTO 0);
    l_sum_qty_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
    l_sum_base_price_cmd_valid : OUT STD_LOGIC;
    l_sum_base_price_cmd_ready : IN STD_LOGIC;
    l_sum_base_price_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
    l_sum_base_price_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
    l_sum_base_price_cmd_ctrl : OUT STD_LOGIC_VECTOR(L_SUM_BASE_PRICE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
    l_sum_base_price_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
    l_sum_disc_price_cmd_valid : OUT STD_LOGIC;
    l_sum_disc_price_cmd_ready : IN STD_LOGIC;
    l_sum_disc_price_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
    l_sum_disc_price_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
    l_sum_disc_price_cmd_ctrl : OUT STD_LOGIC_VECTOR(L_SUM_DISC_PRICE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
    l_sum_disc_price_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
    l_sum_charge_cmd_valid : OUT STD_LOGIC;
    l_sum_charge_cmd_ready : IN STD_LOGIC;
    l_sum_charge_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
    l_sum_charge_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
    l_sum_charge_cmd_ctrl : OUT STD_LOGIC_VECTOR(L_SUM_CHARGE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
    l_sum_charge_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
    l_avg_qty_cmd_valid : OUT STD_LOGIC;
    l_avg_qty_cmd_ready : IN STD_LOGIC;
    l_avg_qty_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
    l_avg_qty_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
    l_avg_qty_cmd_ctrl : OUT STD_LOGIC_VECTOR(L_AVG_QTY_BUS_ADDR_WIDTH - 1 DOWNTO 0);
    l_avg_qty_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
    l_avg_price_cmd_valid : OUT STD_LOGIC;
    l_avg_price_cmd_ready : IN STD_LOGIC;
    l_avg_price_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
    l_avg_price_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
    l_avg_price_cmd_ctrl : OUT STD_LOGIC_VECTOR(L_AVG_PRICE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
    l_avg_price_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
    l_avg_disc_cmd_valid : OUT STD_LOGIC;
    l_avg_disc_cmd_ready : IN STD_LOGIC;
    l_avg_disc_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
    l_avg_disc_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
    l_avg_disc_cmd_ctrl : OUT STD_LOGIC_VECTOR(L_AVG_DISC_BUS_ADDR_WIDTH - 1 DOWNTO 0);
    l_avg_disc_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
    l_count_order_cmd_valid : OUT STD_LOGIC;
    l_count_order_cmd_ready : IN STD_LOGIC;
    l_count_order_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
    l_count_order_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
    l_count_order_cmd_ctrl : OUT STD_LOGIC_VECTOR(L_COUNT_ORDER_BUS_ADDR_WIDTH - 1 DOWNTO 0);
    l_count_order_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0)
  );
END ENTITY;

ARCHITECTURE Implementation OF PriceSummary_Nucleus IS
  COMPONENT PriceSummary IS
    GENERIC (
      INDEX_WIDTH : INTEGER := 32;
      TAG_WIDTH : INTEGER := 1
    );
    PORT (
      kcd_clk : IN STD_LOGIC;
      kcd_reset : IN STD_LOGIC;
      l_quantity_valid : IN STD_LOGIC;
      l_quantity_ready : OUT STD_LOGIC;
      l_quantity_dvalid : IN STD_LOGIC;
      l_quantity_last : IN STD_LOGIC;
      l_quantity : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_extendedprice_valid : IN STD_LOGIC;
      l_extendedprice_ready : OUT STD_LOGIC;
      l_extendedprice_dvalid : IN STD_LOGIC;
      l_extendedprice_last : IN STD_LOGIC;
      l_extendedprice : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_discount_valid : IN STD_LOGIC;
      l_discount_ready : OUT STD_LOGIC;
      l_discount_dvalid : IN STD_LOGIC;
      l_discount_last : IN STD_LOGIC;
      l_discount : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_tax_valid : IN STD_LOGIC;
      l_tax_ready : OUT STD_LOGIC;
      l_tax_dvalid : IN STD_LOGIC;
      l_tax_last : IN STD_LOGIC;
      l_tax : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_returnflag_valid : IN STD_LOGIC;
      l_returnflag_ready : OUT STD_LOGIC;
      l_returnflag_dvalid : IN STD_LOGIC;
      l_returnflag_last : IN STD_LOGIC;
      l_returnflag_length : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      l_returnflag_count : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      l_returnflag_chars_valid : IN STD_LOGIC;
      l_returnflag_chars_ready : OUT STD_LOGIC;
      l_returnflag_chars_dvalid : IN STD_LOGIC;
      l_returnflag_chars_last : IN STD_LOGIC;
      l_returnflag_chars : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      l_returnflag_chars_count : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      l_linestatus_valid : IN STD_LOGIC;
      l_linestatus_ready : OUT STD_LOGIC;
      l_linestatus_dvalid : IN STD_LOGIC;
      l_linestatus_last : IN STD_LOGIC;
      l_linestatus_length : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      l_linestatus_count : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      l_linestatus_chars_valid : IN STD_LOGIC;
      l_linestatus_chars_ready : OUT STD_LOGIC;
      l_linestatus_chars_dvalid : IN STD_LOGIC;
      l_linestatus_chars_last : IN STD_LOGIC;
      l_linestatus_chars : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      l_linestatus_chars_count : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      l_shipdate_valid : IN STD_LOGIC;
      l_shipdate_ready : OUT STD_LOGIC;
      l_shipdate_dvalid : IN STD_LOGIC;
      l_shipdate_last : IN STD_LOGIC;
      l_shipdate : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      l_quantity_unl_valid : IN STD_LOGIC;
      l_quantity_unl_ready : OUT STD_LOGIC;
      l_quantity_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_extendedprice_unl_valid : IN STD_LOGIC;
      l_extendedprice_unl_ready : OUT STD_LOGIC;
      l_extendedprice_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_discount_unl_valid : IN STD_LOGIC;
      l_discount_unl_ready : OUT STD_LOGIC;
      l_discount_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_tax_unl_valid : IN STD_LOGIC;
      l_tax_unl_ready : OUT STD_LOGIC;
      l_tax_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_returnflag_unl_valid : IN STD_LOGIC;
      l_returnflag_unl_ready : OUT STD_LOGIC;
      l_returnflag_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_linestatus_unl_valid : IN STD_LOGIC;
      l_linestatus_unl_ready : OUT STD_LOGIC;
      l_linestatus_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_shipdate_unl_valid : IN STD_LOGIC;
      l_shipdate_unl_ready : OUT STD_LOGIC;
      l_shipdate_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_quantity_cmd_valid : OUT STD_LOGIC;
      l_quantity_cmd_ready : IN STD_LOGIC;
      l_quantity_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_quantity_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_quantity_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_extendedprice_cmd_valid : OUT STD_LOGIC;
      l_extendedprice_cmd_ready : IN STD_LOGIC;
      l_extendedprice_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_extendedprice_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_extendedprice_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_discount_cmd_valid : OUT STD_LOGIC;
      l_discount_cmd_ready : IN STD_LOGIC;
      l_discount_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_discount_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_discount_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_tax_cmd_valid : OUT STD_LOGIC;
      l_tax_cmd_ready : IN STD_LOGIC;
      l_tax_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_tax_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_tax_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_returnflag_cmd_valid : OUT STD_LOGIC;
      l_returnflag_cmd_ready : IN STD_LOGIC;
      l_returnflag_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_returnflag_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_returnflag_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_linestatus_cmd_valid : OUT STD_LOGIC;
      l_linestatus_cmd_ready : IN STD_LOGIC;
      l_linestatus_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_linestatus_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_linestatus_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_shipdate_cmd_valid : OUT STD_LOGIC;
      l_shipdate_cmd_ready : IN STD_LOGIC;
      l_shipdate_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_shipdate_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_shipdate_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_returnflag_o_valid : OUT STD_LOGIC;
      l_returnflag_o_ready : IN STD_LOGIC;
      l_returnflag_o_dvalid : OUT STD_LOGIC;
      l_returnflag_o_last : OUT STD_LOGIC;
      l_returnflag_o_length : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
      l_returnflag_o_count : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      l_returnflag_o_chars_valid : OUT STD_LOGIC;
      l_returnflag_o_chars_ready : IN STD_LOGIC;
      l_returnflag_o_chars_dvalid : OUT STD_LOGIC;
      l_returnflag_o_chars_last : OUT STD_LOGIC;
      l_returnflag_o_chars : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
      l_returnflag_o_chars_count : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      l_linestatus_o_valid : OUT STD_LOGIC;
      l_linestatus_o_ready : IN STD_LOGIC;
      l_linestatus_o_dvalid : OUT STD_LOGIC;
      l_linestatus_o_last : OUT STD_LOGIC;
      l_linestatus_o_length : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
      l_linestatus_o_count : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      l_linestatus_o_chars_valid : OUT STD_LOGIC;
      l_linestatus_o_chars_ready : IN STD_LOGIC;
      l_linestatus_o_chars_dvalid : OUT STD_LOGIC;
      l_linestatus_o_chars_last : OUT STD_LOGIC;
      l_linestatus_o_chars : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
      l_linestatus_o_chars_count : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      l_sum_qty_valid : OUT STD_LOGIC;
      l_sum_qty_ready : IN STD_LOGIC;
      l_sum_qty_dvalid : OUT STD_LOGIC;
      l_sum_qty_last : OUT STD_LOGIC;
      l_sum_qty : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_sum_base_price_valid : OUT STD_LOGIC;
      l_sum_base_price_ready : IN STD_LOGIC;
      l_sum_base_price_dvalid : OUT STD_LOGIC;
      l_sum_base_price_last : OUT STD_LOGIC;
      l_sum_base_price : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_sum_disc_price_valid : OUT STD_LOGIC;
      l_sum_disc_price_ready : IN STD_LOGIC;
      l_sum_disc_price_dvalid : OUT STD_LOGIC;
      l_sum_disc_price_last : OUT STD_LOGIC;
      l_sum_disc_price : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_sum_charge_valid : OUT STD_LOGIC;
      l_sum_charge_ready : IN STD_LOGIC;
      l_sum_charge_dvalid : OUT STD_LOGIC;
      l_sum_charge_last : OUT STD_LOGIC;
      l_sum_charge : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_avg_qty_valid : OUT STD_LOGIC;
      l_avg_qty_ready : IN STD_LOGIC;
      l_avg_qty_dvalid : OUT STD_LOGIC;
      l_avg_qty_last : OUT STD_LOGIC;
      l_avg_qty : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_avg_price_valid : OUT STD_LOGIC;
      l_avg_price_ready : IN STD_LOGIC;
      l_avg_price_dvalid : OUT STD_LOGIC;
      l_avg_price_last : OUT STD_LOGIC;
      l_avg_price : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_avg_disc_valid : OUT STD_LOGIC;
      l_avg_disc_ready : IN STD_LOGIC;
      l_avg_disc_dvalid : OUT STD_LOGIC;
      l_avg_disc_last : OUT STD_LOGIC;
      l_avg_disc : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_count_order_valid : OUT STD_LOGIC;
      l_count_order_ready : IN STD_LOGIC;
      l_count_order_dvalid : OUT STD_LOGIC;
      l_count_order_last : OUT STD_LOGIC;
      l_count_order : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_returnflag_o_unl_valid : IN STD_LOGIC;
      l_returnflag_o_unl_ready : OUT STD_LOGIC;
      l_returnflag_o_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_linestatus_o_unl_valid : IN STD_LOGIC;
      l_linestatus_o_unl_ready : OUT STD_LOGIC;
      l_linestatus_o_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_sum_qty_unl_valid : IN STD_LOGIC;
      l_sum_qty_unl_ready : OUT STD_LOGIC;
      l_sum_qty_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_sum_base_price_unl_valid : IN STD_LOGIC;
      l_sum_base_price_unl_ready : OUT STD_LOGIC;
      l_sum_base_price_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_sum_disc_price_unl_valid : IN STD_LOGIC;
      l_sum_disc_price_unl_ready : OUT STD_LOGIC;
      l_sum_disc_price_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_sum_charge_unl_valid : IN STD_LOGIC;
      l_sum_charge_unl_ready : OUT STD_LOGIC;
      l_sum_charge_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_avg_qty_unl_valid : IN STD_LOGIC;
      l_avg_qty_unl_ready : OUT STD_LOGIC;
      l_avg_qty_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_avg_price_unl_valid : IN STD_LOGIC;
      l_avg_price_unl_ready : OUT STD_LOGIC;
      l_avg_price_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_avg_disc_unl_valid : IN STD_LOGIC;
      l_avg_disc_unl_ready : OUT STD_LOGIC;
      l_avg_disc_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_count_order_unl_valid : IN STD_LOGIC;
      l_count_order_unl_ready : OUT STD_LOGIC;
      l_count_order_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_returnflag_o_cmd_valid : OUT STD_LOGIC;
      l_returnflag_o_cmd_ready : IN STD_LOGIC;
      l_returnflag_o_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_returnflag_o_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_returnflag_o_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_linestatus_o_cmd_valid : OUT STD_LOGIC;
      l_linestatus_o_cmd_ready : IN STD_LOGIC;
      l_linestatus_o_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_linestatus_o_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_linestatus_o_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_sum_qty_cmd_valid : OUT STD_LOGIC;
      l_sum_qty_cmd_ready : IN STD_LOGIC;
      l_sum_qty_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_sum_qty_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_sum_qty_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_sum_base_price_cmd_valid : OUT STD_LOGIC;
      l_sum_base_price_cmd_ready : IN STD_LOGIC;
      l_sum_base_price_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_sum_base_price_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_sum_base_price_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_sum_disc_price_cmd_valid : OUT STD_LOGIC;
      l_sum_disc_price_cmd_ready : IN STD_LOGIC;
      l_sum_disc_price_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_sum_disc_price_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_sum_disc_price_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_sum_charge_cmd_valid : OUT STD_LOGIC;
      l_sum_charge_cmd_ready : IN STD_LOGIC;
      l_sum_charge_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_sum_charge_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_sum_charge_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_avg_qty_cmd_valid : OUT STD_LOGIC;
      l_avg_qty_cmd_ready : IN STD_LOGIC;
      l_avg_qty_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_avg_qty_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_avg_qty_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_avg_price_cmd_valid : OUT STD_LOGIC;
      l_avg_price_cmd_ready : IN STD_LOGIC;
      l_avg_price_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_avg_price_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_avg_price_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_avg_disc_cmd_valid : OUT STD_LOGIC;
      l_avg_disc_cmd_ready : IN STD_LOGIC;
      l_avg_disc_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_avg_disc_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_avg_disc_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_count_order_cmd_valid : OUT STD_LOGIC;
      l_count_order_cmd_ready : IN STD_LOGIC;
      l_count_order_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_count_order_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_count_order_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      start : IN STD_LOGIC;
      stop : IN STD_LOGIC;
      reset : IN STD_LOGIC;
      idle : OUT STD_LOGIC;
      busy : OUT STD_LOGIC;
      done : OUT STD_LOGIC;
      result : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_firstidx : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      l_lastidx : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      rhigh : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
      rlow : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
      status_1 : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
      status_2 : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
      r1 : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
      r2 : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
      r3 : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
      r4 : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
      r5 : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
      r6 : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
      r7 : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
      r8 : OUT STD_LOGIC_VECTOR(63 DOWNTO 0)
    );
  END COMPONENT;

  SIGNAL PriceSummary_inst_l_quantity_valid : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_quantity_ready : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_quantity_dvalid : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_quantity_last : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_quantity : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummary_inst_l_extendedprice_valid : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_extendedprice_ready : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_extendedprice_dvalid : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_extendedprice_last : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_extendedprice : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummary_inst_l_discount_valid : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_discount_ready : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_discount_dvalid : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_discount_last : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_discount : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummary_inst_l_tax_valid : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_tax_ready : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_tax_dvalid : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_tax_last : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_tax : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummary_inst_l_returnflag_valid : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_returnflag_ready : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_returnflag_dvalid : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_returnflag_last : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_returnflag_length : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummary_inst_l_returnflag_count : STD_LOGIC_VECTOR(0 DOWNTO 0);
  SIGNAL PriceSummary_inst_l_returnflag_chars_valid : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_returnflag_chars_ready : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_returnflag_chars_dvalid : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_returnflag_chars_last : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_returnflag_chars : STD_LOGIC_VECTOR(7 DOWNTO 0);
  SIGNAL PriceSummary_inst_l_returnflag_chars_count : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummary_inst_l_linestatus_valid : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_linestatus_ready : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_linestatus_dvalid : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_linestatus_last : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_linestatus_length : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummary_inst_l_linestatus_count : STD_LOGIC_VECTOR(0 DOWNTO 0);
  SIGNAL PriceSummary_inst_l_linestatus_chars_valid : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_linestatus_chars_ready : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_linestatus_chars_dvalid : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_linestatus_chars_last : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_linestatus_chars : STD_LOGIC_VECTOR(7 DOWNTO 0);
  SIGNAL PriceSummary_inst_l_linestatus_chars_count : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummary_inst_l_shipdate_valid : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_shipdate_ready : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_shipdate_dvalid : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_shipdate_last : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_shipdate : STD_LOGIC_VECTOR(31 DOWNTO 0);

  SIGNAL PriceSummary_inst_l_quantity_unl_valid : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_quantity_unl_ready : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_quantity_unl_tag : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummary_inst_l_extendedprice_unl_valid : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_extendedprice_unl_ready : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_extendedprice_unl_tag : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummary_inst_l_discount_unl_valid : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_discount_unl_ready : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_discount_unl_tag : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummary_inst_l_tax_unl_valid : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_tax_unl_ready : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_tax_unl_tag : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummary_inst_l_returnflag_unl_valid : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_returnflag_unl_ready : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_returnflag_unl_tag : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummary_inst_l_linestatus_unl_valid : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_linestatus_unl_ready : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_linestatus_unl_tag : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummary_inst_l_shipdate_unl_valid : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_shipdate_unl_ready : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_shipdate_unl_tag : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummary_inst_l_quantity_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_quantity_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_quantity_cmd_firstIdx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummary_inst_l_quantity_cmd_lastIdx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummary_inst_l_quantity_cmd_tag : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummary_inst_l_extendedprice_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_extendedprice_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_extendedprice_cmd_firstIdx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummary_inst_l_extendedprice_cmd_lastIdx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummary_inst_l_extendedprice_cmd_tag : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummary_inst_l_discount_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_discount_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_discount_cmd_firstIdx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummary_inst_l_discount_cmd_lastIdx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummary_inst_l_discount_cmd_tag : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummary_inst_l_tax_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_tax_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_tax_cmd_firstIdx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummary_inst_l_tax_cmd_lastIdx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummary_inst_l_tax_cmd_tag : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummary_inst_l_returnflag_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_returnflag_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_returnflag_cmd_firstIdx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummary_inst_l_returnflag_cmd_lastIdx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummary_inst_l_returnflag_cmd_tag : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummary_inst_l_linestatus_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_linestatus_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_linestatus_cmd_firstIdx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummary_inst_l_linestatus_cmd_lastIdx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummary_inst_l_linestatus_cmd_tag : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummary_inst_l_shipdate_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_shipdate_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummary_inst_l_shipdate_cmd_firstIdx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummary_inst_l_shipdate_cmd_lastIdx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummary_inst_l_shipdate_cmd_tag : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummaryWriter_inst_l_returnflag_o_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_returnflag_o_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_returnflag_o_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_returnflag_o_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_returnflag_o_length : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummaryWriter_inst_l_returnflag_o_count : STD_LOGIC_VECTOR(0 DOWNTO 0);
  SIGNAL PriceSummaryWriter_inst_l_returnflag_o_chars_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_returnflag_o_chars_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_returnflag_o_chars_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_returnflag_o_chars_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_returnflag_o_chars : STD_LOGIC_VECTOR(7 DOWNTO 0);
  SIGNAL PriceSummaryWriter_inst_l_returnflag_o_chars_count : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummaryWriter_inst_l_linestatus_o_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_linestatus_o_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_linestatus_o_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_linestatus_o_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_linestatus_o_length : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummaryWriter_inst_l_linestatus_o_count : STD_LOGIC_VECTOR(0 DOWNTO 0);
  SIGNAL PriceSummaryWriter_inst_l_linestatus_o_chars_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_linestatus_o_chars_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_linestatus_o_chars_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_linestatus_o_chars_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_linestatus_o_chars : STD_LOGIC_VECTOR(7 DOWNTO 0);
  SIGNAL PriceSummaryWriter_inst_l_linestatus_o_chars_count : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummaryWriter_inst_l_sum_qty_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_sum_qty_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_sum_qty_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_sum_qty_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_sum_qty : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummaryWriter_inst_l_sum_base_price_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_sum_base_price_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_sum_base_price_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_sum_base_price_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_sum_base_price : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummaryWriter_inst_l_sum_disc_price_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_sum_disc_price_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_sum_disc_price_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_sum_disc_price_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_sum_disc_price : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummaryWriter_inst_l_sum_charge_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_sum_charge_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_sum_charge_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_sum_charge_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_sum_charge : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummaryWriter_inst_l_avg_qty_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_avg_qty_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_avg_qty_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_avg_qty_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_avg_qty : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummaryWriter_inst_l_avg_price_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_avg_price_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_avg_price_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_avg_price_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_avg_price : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummaryWriter_inst_l_avg_disc_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_avg_disc_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_avg_disc_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_avg_disc_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_avg_disc : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummaryWriter_inst_l_count_order_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_count_order_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_count_order_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_count_order_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_count_order : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummaryWriter_inst_l_returnflag_o_unl_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_returnflag_o_unl_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_returnflag_o_unl_tag : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummaryWriter_inst_l_linestatus_o_unl_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_linestatus_o_unl_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_linestatus_o_unl_tag : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummaryWriter_inst_l_sum_qty_unl_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_sum_qty_unl_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_sum_qty_unl_tag : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummaryWriter_inst_l_sum_base_price_unl_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_sum_base_price_unl_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_sum_base_price_unl_tag : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummaryWriter_inst_l_sum_disc_price_unl_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_sum_disc_price_unl_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_sum_disc_price_unl_tag : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummaryWriter_inst_l_sum_charge_unl_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_sum_charge_unl_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_sum_charge_unl_tag : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummaryWriter_inst_l_avg_qty_unl_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_avg_qty_unl_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_avg_qty_unl_tag : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummaryWriter_inst_l_avg_price_unl_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_avg_price_unl_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_avg_price_unl_tag : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummaryWriter_inst_l_avg_disc_unl_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_avg_disc_unl_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_avg_disc_unl_tag : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummaryWriter_inst_l_count_order_unl_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_count_order_unl_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_count_order_unl_tag : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummaryWriter_inst_l_returnflag_o_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_returnflag_o_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_returnflag_o_cmd_firstIdx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummaryWriter_inst_l_returnflag_o_cmd_lastIdx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummaryWriter_inst_l_returnflag_o_cmd_tag : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummaryWriter_inst_l_linestatus_o_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_linestatus_o_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_linestatus_o_cmd_firstIdx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummaryWriter_inst_l_linestatus_o_cmd_lastIdx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummaryWriter_inst_l_linestatus_o_cmd_tag : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummaryWriter_inst_l_sum_qty_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_sum_qty_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_sum_qty_cmd_firstIdx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummaryWriter_inst_l_sum_qty_cmd_lastIdx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummaryWriter_inst_l_sum_qty_cmd_tag : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummaryWriter_inst_l_sum_base_price_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_sum_base_price_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_sum_base_price_cmd_firstIdx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummaryWriter_inst_l_sum_base_price_cmd_lastIdx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummaryWriter_inst_l_sum_base_price_cmd_tag : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummaryWriter_inst_l_sum_disc_price_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_sum_disc_price_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_sum_disc_price_cmd_firstIdx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummaryWriter_inst_l_sum_disc_price_cmd_lastIdx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummaryWriter_inst_l_sum_disc_price_cmd_tag : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummaryWriter_inst_l_sum_charge_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_sum_charge_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_sum_charge_cmd_firstIdx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummaryWriter_inst_l_sum_charge_cmd_lastIdx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummaryWriter_inst_l_sum_charge_cmd_tag : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummaryWriter_inst_l_avg_qty_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_avg_qty_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_avg_qty_cmd_firstIdx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummaryWriter_inst_l_avg_qty_cmd_lastIdx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummaryWriter_inst_l_avg_qty_cmd_tag : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummaryWriter_inst_l_avg_price_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_avg_price_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_avg_price_cmd_firstIdx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummaryWriter_inst_l_avg_price_cmd_lastIdx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummaryWriter_inst_l_avg_price_cmd_tag : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummaryWriter_inst_l_avg_disc_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_avg_disc_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_avg_disc_cmd_firstIdx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummaryWriter_inst_l_avg_disc_cmd_lastIdx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummaryWriter_inst_l_avg_disc_cmd_tag : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummaryWriter_inst_l_count_order_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_count_order_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_inst_l_count_order_cmd_firstIdx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummaryWriter_inst_l_count_order_cmd_lastIdx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummaryWriter_inst_l_count_order_cmd_tag : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummary_inst_start : STD_LOGIC;
  SIGNAL PriceSummary_inst_stop : STD_LOGIC;
  SIGNAL PriceSummary_inst_reset : STD_LOGIC;
  SIGNAL PriceSummary_inst_idle : STD_LOGIC;
  SIGNAL PriceSummary_inst_busy : STD_LOGIC;
  SIGNAL PriceSummary_inst_done : STD_LOGIC;
  SIGNAL PriceSummary_inst_result : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL PriceSummary_inst_l_firstidx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummary_inst_l_lastidx : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummary_inst_rhigh : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummary_inst_rlow : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummary_inst_status_1 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummary_inst_status_2 : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummary_inst_r1 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL PriceSummary_inst_r2 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL PriceSummary_inst_r3 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL PriceSummary_inst_r4 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL PriceSummary_inst_r5 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL PriceSummary_inst_r6 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL PriceSummary_inst_r7 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL PriceSummary_inst_r8 : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL mmio_inst_f_start_data : STD_LOGIC;
  SIGNAL mmio_inst_f_stop_data : STD_LOGIC;
  SIGNAL mmio_inst_f_reset_data : STD_LOGIC;
  SIGNAL mmio_inst_f_idle_write_data : STD_LOGIC;
  SIGNAL mmio_inst_f_busy_write_data : STD_LOGIC;
  SIGNAL mmio_inst_f_done_write_data : STD_LOGIC;
  SIGNAL mmio_inst_f_result_write_data : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL mmio_inst_f_l_firstidx_data : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL mmio_inst_f_l_lastidx_data : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL mmio_inst_f_l_quantity_values_data : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL mmio_inst_f_l_extendedprice_values_data : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL mmio_inst_f_l_discount_values_data : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL mmio_inst_f_l_tax_values_data : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL mmio_inst_f_l_returnflag_offsets_data : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL mmio_inst_f_l_returnflag_values_data : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL mmio_inst_f_l_linestatus_offsets_data : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL mmio_inst_f_l_linestatus_values_data : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL mmio_inst_f_l_shipdate_values_data : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL mmio_inst_f_l_returnflag_o_offsets_data : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL mmio_inst_f_l_returnflag_o_values_data : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL mmio_inst_f_l_linestatus_o_offsets_data : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL mmio_inst_f_l_linestatus_o_values_data : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL mmio_inst_f_l_sum_qty_values_data : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL mmio_inst_f_l_sum_base_price_values_data : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL mmio_inst_f_l_sum_disc_price_values_data : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL mmio_inst_f_l_sum_charge_values_data : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL mmio_inst_f_l_avg_qty_values_data : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL mmio_inst_f_l_avg_price_values_data : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL mmio_inst_f_l_avg_disc_values_data : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL mmio_inst_f_l_count_order_values_data : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL mmio_inst_f_rhigh_write_data : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL mmio_inst_f_rlow_write_data : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL mmio_inst_f_status_1_write_data : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL mmio_inst_f_status_2_write_data : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL mmio_inst_f_r1_write_data : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL mmio_inst_f_r2_write_data : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL mmio_inst_f_r3_write_data : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL mmio_inst_f_r4_write_data : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL mmio_inst_f_r5_write_data : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL mmio_inst_f_r6_write_data : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL mmio_inst_f_r7_write_data : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL mmio_inst_f_r8_write_data : STD_LOGIC_VECTOR(63 DOWNTO 0);
  SIGNAL mmio_inst_f_Profile_enable_data : STD_LOGIC;
  SIGNAL mmio_inst_f_Profile_clear_data : STD_LOGIC;
  SIGNAL mmio_inst_mmio_awvalid : STD_LOGIC;
  SIGNAL mmio_inst_mmio_awready : STD_LOGIC;
  SIGNAL mmio_inst_mmio_awaddr : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL mmio_inst_mmio_wvalid : STD_LOGIC;
  SIGNAL mmio_inst_mmio_wready : STD_LOGIC;
  SIGNAL mmio_inst_mmio_wdata : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL mmio_inst_mmio_wstrb : STD_LOGIC_VECTOR(3 DOWNTO 0);
  SIGNAL mmio_inst_mmio_bvalid : STD_LOGIC;
  SIGNAL mmio_inst_mmio_bready : STD_LOGIC;
  SIGNAL mmio_inst_mmio_bresp : STD_LOGIC_VECTOR(1 DOWNTO 0);
  SIGNAL mmio_inst_mmio_arvalid : STD_LOGIC;
  SIGNAL mmio_inst_mmio_arready : STD_LOGIC;
  SIGNAL mmio_inst_mmio_araddr : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL mmio_inst_mmio_rvalid : STD_LOGIC;
  SIGNAL mmio_inst_mmio_rready : STD_LOGIC;
  SIGNAL mmio_inst_mmio_rdata : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL mmio_inst_mmio_rresp : STD_LOGIC_VECTOR(1 DOWNTO 0);

  SIGNAL l_quantity_cmd_accm_inst_kernel_cmd_valid : STD_LOGIC;
  SIGNAL l_quantity_cmd_accm_inst_kernel_cmd_ready : STD_LOGIC;
  SIGNAL l_quantity_cmd_accm_inst_kernel_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_quantity_cmd_accm_inst_kernel_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_quantity_cmd_accm_inst_kernel_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL l_quantity_cmd_accm_inst_nucleus_cmd_valid : STD_LOGIC;
  SIGNAL l_quantity_cmd_accm_inst_nucleus_cmd_ready : STD_LOGIC;
  SIGNAL l_quantity_cmd_accm_inst_nucleus_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_quantity_cmd_accm_inst_nucleus_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_quantity_cmd_accm_inst_nucleus_cmd_ctrl : STD_LOGIC_VECTOR(L_QUANTITY_BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL l_quantity_cmd_accm_inst_nucleus_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL l_extendedprice_cmd_accm_inst_kernel_cmd_valid : STD_LOGIC;
  SIGNAL l_extendedprice_cmd_accm_inst_kernel_cmd_ready : STD_LOGIC;
  SIGNAL l_extendedprice_cmd_accm_inst_kernel_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_extendedprice_cmd_accm_inst_kernel_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_extendedprice_cmd_accm_inst_kernel_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL l_extendedprice_cmd_accm_inst_nucleus_cmd_valid : STD_LOGIC;
  SIGNAL l_extendedprice_cmd_accm_inst_nucleus_cmd_ready : STD_LOGIC;
  SIGNAL l_extendedprice_cmd_accm_inst_nucleus_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_extendedprice_cmd_accm_inst_nucleus_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_extendedprice_cmd_accm_inst_nucleus_cmd_ctrl : STD_LOGIC_VECTOR(L_EXTENDEDPRICE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL l_extendedprice_cmd_accm_inst_nucleus_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL l_discount_cmd_accm_inst_kernel_cmd_valid : STD_LOGIC;
  SIGNAL l_discount_cmd_accm_inst_kernel_cmd_ready : STD_LOGIC;
  SIGNAL l_discount_cmd_accm_inst_kernel_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_discount_cmd_accm_inst_kernel_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_discount_cmd_accm_inst_kernel_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL l_discount_cmd_accm_inst_nucleus_cmd_valid : STD_LOGIC;
  SIGNAL l_discount_cmd_accm_inst_nucleus_cmd_ready : STD_LOGIC;
  SIGNAL l_discount_cmd_accm_inst_nucleus_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_discount_cmd_accm_inst_nucleus_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_discount_cmd_accm_inst_nucleus_cmd_ctrl : STD_LOGIC_VECTOR(L_DISCOUNT_BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL l_discount_cmd_accm_inst_nucleus_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL l_tax_cmd_accm_inst_kernel_cmd_valid : STD_LOGIC;
  SIGNAL l_tax_cmd_accm_inst_kernel_cmd_ready : STD_LOGIC;
  SIGNAL l_tax_cmd_accm_inst_kernel_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_tax_cmd_accm_inst_kernel_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_tax_cmd_accm_inst_kernel_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL l_tax_cmd_accm_inst_nucleus_cmd_valid : STD_LOGIC;
  SIGNAL l_tax_cmd_accm_inst_nucleus_cmd_ready : STD_LOGIC;
  SIGNAL l_tax_cmd_accm_inst_nucleus_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_tax_cmd_accm_inst_nucleus_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_tax_cmd_accm_inst_nucleus_cmd_ctrl : STD_LOGIC_VECTOR(L_TAX_BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL l_tax_cmd_accm_inst_nucleus_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL l_returnflag_cmd_accm_inst_kernel_cmd_valid : STD_LOGIC;
  SIGNAL l_returnflag_cmd_accm_inst_kernel_cmd_ready : STD_LOGIC;
  SIGNAL l_returnflag_cmd_accm_inst_kernel_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_returnflag_cmd_accm_inst_kernel_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_returnflag_cmd_accm_inst_kernel_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL l_returnflag_cmd_accm_inst_nucleus_cmd_valid : STD_LOGIC;
  SIGNAL l_returnflag_cmd_accm_inst_nucleus_cmd_ready : STD_LOGIC;
  SIGNAL l_returnflag_cmd_accm_inst_nucleus_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_returnflag_cmd_accm_inst_nucleus_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_returnflag_cmd_accm_inst_nucleus_cmd_ctrl : STD_LOGIC_VECTOR(2 * L_RETURNFLAG_BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL l_returnflag_cmd_accm_inst_nucleus_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL l_linestatus_cmd_accm_inst_kernel_cmd_valid : STD_LOGIC;
  SIGNAL l_linestatus_cmd_accm_inst_kernel_cmd_ready : STD_LOGIC;
  SIGNAL l_linestatus_cmd_accm_inst_kernel_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_linestatus_cmd_accm_inst_kernel_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_linestatus_cmd_accm_inst_kernel_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL l_linestatus_cmd_accm_inst_nucleus_cmd_valid : STD_LOGIC;
  SIGNAL l_linestatus_cmd_accm_inst_nucleus_cmd_ready : STD_LOGIC;
  SIGNAL l_linestatus_cmd_accm_inst_nucleus_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_linestatus_cmd_accm_inst_nucleus_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_linestatus_cmd_accm_inst_nucleus_cmd_ctrl : STD_LOGIC_VECTOR(2 * L_LINESTATUS_BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL l_linestatus_cmd_accm_inst_nucleus_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL l_shipdate_cmd_accm_inst_kernel_cmd_valid : STD_LOGIC;
  SIGNAL l_shipdate_cmd_accm_inst_kernel_cmd_ready : STD_LOGIC;
  SIGNAL l_shipdate_cmd_accm_inst_kernel_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_shipdate_cmd_accm_inst_kernel_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_shipdate_cmd_accm_inst_kernel_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL l_shipdate_cmd_accm_inst_nucleus_cmd_valid : STD_LOGIC;
  SIGNAL l_shipdate_cmd_accm_inst_nucleus_cmd_ready : STD_LOGIC;
  SIGNAL l_shipdate_cmd_accm_inst_nucleus_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_shipdate_cmd_accm_inst_nucleus_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_shipdate_cmd_accm_inst_nucleus_cmd_ctrl : STD_LOGIC_VECTOR(L_SHIPDATE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL l_shipdate_cmd_accm_inst_nucleus_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL l_quantity_cmd_accm_inst_ctrl : STD_LOGIC_VECTOR(L_QUANTITY_BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL l_extendedprice_cmd_accm_inst_ctrl : STD_LOGIC_VECTOR(L_EXTENDEDPRICE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL l_discount_cmd_accm_inst_ctrl : STD_LOGIC_VECTOR(L_DISCOUNT_BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL l_tax_cmd_accm_inst_ctrl : STD_LOGIC_VECTOR(L_TAX_BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL l_returnflag_cmd_accm_inst_ctrl : STD_LOGIC_VECTOR(2 * L_RETURNFLAG_BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL l_linestatus_cmd_accm_inst_ctrl : STD_LOGIC_VECTOR(2 * L_LINESTATUS_BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL l_shipdate_cmd_accm_inst_ctrl : STD_LOGIC_VECTOR(L_SHIPDATE_BUS_ADDR_WIDTH - 1 DOWNTO 0);

  SIGNAL l_returnflag_o_cmd_accm_inst_kernel_cmd_valid : STD_LOGIC;
  SIGNAL l_returnflag_o_cmd_accm_inst_kernel_cmd_ready : STD_LOGIC;
  SIGNAL l_returnflag_o_cmd_accm_inst_kernel_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_returnflag_o_cmd_accm_inst_kernel_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_returnflag_o_cmd_accm_inst_kernel_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL l_returnflag_o_cmd_accm_inst_nucleus_cmd_valid : STD_LOGIC;
  SIGNAL l_returnflag_o_cmd_accm_inst_nucleus_cmd_ready : STD_LOGIC;
  SIGNAL l_returnflag_o_cmd_accm_inst_nucleus_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_returnflag_o_cmd_accm_inst_nucleus_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_returnflag_o_cmd_accm_inst_nucleus_cmd_ctrl : STD_LOGIC_VECTOR(2 * L_RETURNFLAG_O_BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL l_returnflag_o_cmd_accm_inst_nucleus_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL l_linestatus_o_cmd_accm_inst_kernel_cmd_valid : STD_LOGIC;
  SIGNAL l_linestatus_o_cmd_accm_inst_kernel_cmd_ready : STD_LOGIC;
  SIGNAL l_linestatus_o_cmd_accm_inst_kernel_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_linestatus_o_cmd_accm_inst_kernel_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_linestatus_o_cmd_accm_inst_kernel_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL l_linestatus_o_cmd_accm_inst_nucleus_cmd_valid : STD_LOGIC;
  SIGNAL l_linestatus_o_cmd_accm_inst_nucleus_cmd_ready : STD_LOGIC;
  SIGNAL l_linestatus_o_cmd_accm_inst_nucleus_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_linestatus_o_cmd_accm_inst_nucleus_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_linestatus_o_cmd_accm_inst_nucleus_cmd_ctrl : STD_LOGIC_VECTOR(2 * L_LINESTATUS_O_BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL l_linestatus_o_cmd_accm_inst_nucleus_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL l_sum_qty_cmd_accm_inst_kernel_cmd_valid : STD_LOGIC;
  SIGNAL l_sum_qty_cmd_accm_inst_kernel_cmd_ready : STD_LOGIC;
  SIGNAL l_sum_qty_cmd_accm_inst_kernel_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_sum_qty_cmd_accm_inst_kernel_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_sum_qty_cmd_accm_inst_kernel_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL l_sum_qty_cmd_accm_inst_nucleus_cmd_valid : STD_LOGIC;
  SIGNAL l_sum_qty_cmd_accm_inst_nucleus_cmd_ready : STD_LOGIC;
  SIGNAL l_sum_qty_cmd_accm_inst_nucleus_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_sum_qty_cmd_accm_inst_nucleus_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_sum_qty_cmd_accm_inst_nucleus_cmd_ctrl : STD_LOGIC_VECTOR(L_SUM_QTY_BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL l_sum_qty_cmd_accm_inst_nucleus_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL l_sum_base_price_cmd_accm_inst_kernel_cmd_valid : STD_LOGIC;
  SIGNAL l_sum_base_price_cmd_accm_inst_kernel_cmd_ready : STD_LOGIC;
  SIGNAL l_sum_base_price_cmd_accm_inst_kernel_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_sum_base_price_cmd_accm_inst_kernel_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_sum_base_price_cmd_accm_inst_kernel_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL l_sum_base_price_cmd_accm_inst_nucleus_cmd_valid : STD_LOGIC;
  SIGNAL l_sum_base_price_cmd_accm_inst_nucleus_cmd_ready : STD_LOGIC;
  SIGNAL l_sum_base_price_cmd_accm_inst_nucleus_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_sum_base_price_cmd_accm_inst_nucleus_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_sum_base_price_cmd_accm_inst_nucleus_cmd_ctrl : STD_LOGIC_VECTOR(L_SUM_BASE_PRICE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL l_sum_base_price_cmd_accm_inst_nucleus_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL l_sum_disc_price_cmd_accm_inst_kernel_cmd_valid : STD_LOGIC;
  SIGNAL l_sum_disc_price_cmd_accm_inst_kernel_cmd_ready : STD_LOGIC;
  SIGNAL l_sum_disc_price_cmd_accm_inst_kernel_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_sum_disc_price_cmd_accm_inst_kernel_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_sum_disc_price_cmd_accm_inst_kernel_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL l_sum_disc_price_cmd_accm_inst_nucleus_cmd_valid : STD_LOGIC;
  SIGNAL l_sum_disc_price_cmd_accm_inst_nucleus_cmd_ready : STD_LOGIC;
  SIGNAL l_sum_disc_price_cmd_accm_inst_nucleus_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_sum_disc_price_cmd_accm_inst_nucleus_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_sum_disc_price_cmd_accm_inst_nucleus_cmd_ctrl : STD_LOGIC_VECTOR(L_SUM_DISC_PRICE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL l_sum_disc_price_cmd_accm_inst_nucleus_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL l_sum_charge_cmd_accm_inst_kernel_cmd_valid : STD_LOGIC;
  SIGNAL l_sum_charge_cmd_accm_inst_kernel_cmd_ready : STD_LOGIC;
  SIGNAL l_sum_charge_cmd_accm_inst_kernel_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_sum_charge_cmd_accm_inst_kernel_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_sum_charge_cmd_accm_inst_kernel_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL l_sum_charge_cmd_accm_inst_nucleus_cmd_valid : STD_LOGIC;
  SIGNAL l_sum_charge_cmd_accm_inst_nucleus_cmd_ready : STD_LOGIC;
  SIGNAL l_sum_charge_cmd_accm_inst_nucleus_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_sum_charge_cmd_accm_inst_nucleus_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_sum_charge_cmd_accm_inst_nucleus_cmd_ctrl : STD_LOGIC_VECTOR(L_SUM_CHARGE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL l_sum_charge_cmd_accm_inst_nucleus_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL l_avg_qty_cmd_accm_inst_kernel_cmd_valid : STD_LOGIC;
  SIGNAL l_avg_qty_cmd_accm_inst_kernel_cmd_ready : STD_LOGIC;
  SIGNAL l_avg_qty_cmd_accm_inst_kernel_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_avg_qty_cmd_accm_inst_kernel_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_avg_qty_cmd_accm_inst_kernel_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL l_avg_qty_cmd_accm_inst_nucleus_cmd_valid : STD_LOGIC;
  SIGNAL l_avg_qty_cmd_accm_inst_nucleus_cmd_ready : STD_LOGIC;
  SIGNAL l_avg_qty_cmd_accm_inst_nucleus_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_avg_qty_cmd_accm_inst_nucleus_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_avg_qty_cmd_accm_inst_nucleus_cmd_ctrl : STD_LOGIC_VECTOR(L_AVG_QTY_BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL l_avg_qty_cmd_accm_inst_nucleus_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL l_avg_price_cmd_accm_inst_kernel_cmd_valid : STD_LOGIC;
  SIGNAL l_avg_price_cmd_accm_inst_kernel_cmd_ready : STD_LOGIC;
  SIGNAL l_avg_price_cmd_accm_inst_kernel_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_avg_price_cmd_accm_inst_kernel_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_avg_price_cmd_accm_inst_kernel_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL l_avg_price_cmd_accm_inst_nucleus_cmd_valid : STD_LOGIC;
  SIGNAL l_avg_price_cmd_accm_inst_nucleus_cmd_ready : STD_LOGIC;
  SIGNAL l_avg_price_cmd_accm_inst_nucleus_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_avg_price_cmd_accm_inst_nucleus_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_avg_price_cmd_accm_inst_nucleus_cmd_ctrl : STD_LOGIC_VECTOR(L_AVG_PRICE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL l_avg_price_cmd_accm_inst_nucleus_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL l_avg_disc_cmd_accm_inst_kernel_cmd_valid : STD_LOGIC;
  SIGNAL l_avg_disc_cmd_accm_inst_kernel_cmd_ready : STD_LOGIC;
  SIGNAL l_avg_disc_cmd_accm_inst_kernel_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_avg_disc_cmd_accm_inst_kernel_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_avg_disc_cmd_accm_inst_kernel_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL l_avg_disc_cmd_accm_inst_nucleus_cmd_valid : STD_LOGIC;
  SIGNAL l_avg_disc_cmd_accm_inst_nucleus_cmd_ready : STD_LOGIC;
  SIGNAL l_avg_disc_cmd_accm_inst_nucleus_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_avg_disc_cmd_accm_inst_nucleus_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_avg_disc_cmd_accm_inst_nucleus_cmd_ctrl : STD_LOGIC_VECTOR(L_AVG_DISC_BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL l_avg_disc_cmd_accm_inst_nucleus_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL l_count_order_cmd_accm_inst_kernel_cmd_valid : STD_LOGIC;
  SIGNAL l_count_order_cmd_accm_inst_kernel_cmd_ready : STD_LOGIC;
  SIGNAL l_count_order_cmd_accm_inst_kernel_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_count_order_cmd_accm_inst_kernel_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_count_order_cmd_accm_inst_kernel_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL l_count_order_cmd_accm_inst_nucleus_cmd_valid : STD_LOGIC;
  SIGNAL l_count_order_cmd_accm_inst_nucleus_cmd_ready : STD_LOGIC;
  SIGNAL l_count_order_cmd_accm_inst_nucleus_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_count_order_cmd_accm_inst_nucleus_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL l_count_order_cmd_accm_inst_nucleus_cmd_ctrl : STD_LOGIC_VECTOR(L_COUNT_ORDER_BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL l_count_order_cmd_accm_inst_nucleus_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL l_returnflag_o_cmd_accm_inst_ctrl : STD_LOGIC_VECTOR(2 * L_RETURNFLAG_O_BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL l_linestatus_o_cmd_accm_inst_ctrl : STD_LOGIC_VECTOR(2 * L_LINESTATUS_O_BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL l_sum_qty_cmd_accm_inst_ctrl : STD_LOGIC_VECTOR(L_SUM_QTY_BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL l_sum_base_price_cmd_accm_inst_ctrl : STD_LOGIC_VECTOR(L_SUM_BASE_PRICE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL l_sum_disc_price_cmd_accm_inst_ctrl : STD_LOGIC_VECTOR(L_SUM_DISC_PRICE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL l_sum_charge_cmd_accm_inst_ctrl : STD_LOGIC_VECTOR(L_SUM_CHARGE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL l_avg_qty_cmd_accm_inst_ctrl : STD_LOGIC_VECTOR(L_AVG_QTY_BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL l_avg_price_cmd_accm_inst_ctrl : STD_LOGIC_VECTOR(L_AVG_PRICE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL l_avg_disc_cmd_accm_inst_ctrl : STD_LOGIC_VECTOR(L_AVG_DISC_BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL l_count_order_cmd_accm_inst_ctrl : STD_LOGIC_VECTOR(L_COUNT_ORDER_BUS_ADDR_WIDTH - 1 DOWNTO 0);
BEGIN
  PriceSummary_inst : PriceSummary
  GENERIC MAP(
    INDEX_WIDTH => 32,
    TAG_WIDTH => 1
  )
  PORT MAP(
    kcd_clk => kcd_clk,
    kcd_reset => kcd_reset,
    l_quantity_valid => PriceSummary_inst_l_quantity_valid,
    l_quantity_ready => PriceSummary_inst_l_quantity_ready,
    l_quantity_dvalid => PriceSummary_inst_l_quantity_dvalid,
    l_quantity_last => PriceSummary_inst_l_quantity_last,
    l_quantity => PriceSummary_inst_l_quantity,
    l_extendedprice_valid => PriceSummary_inst_l_extendedprice_valid,
    l_extendedprice_ready => PriceSummary_inst_l_extendedprice_ready,
    l_extendedprice_dvalid => PriceSummary_inst_l_extendedprice_dvalid,
    l_extendedprice_last => PriceSummary_inst_l_extendedprice_last,
    l_extendedprice => PriceSummary_inst_l_extendedprice,
    l_discount_valid => PriceSummary_inst_l_discount_valid,
    l_discount_ready => PriceSummary_inst_l_discount_ready,
    l_discount_dvalid => PriceSummary_inst_l_discount_dvalid,
    l_discount_last => PriceSummary_inst_l_discount_last,
    l_discount => PriceSummary_inst_l_discount,
    l_tax_valid => PriceSummary_inst_l_tax_valid,
    l_tax_ready => PriceSummary_inst_l_tax_ready,
    l_tax_dvalid => PriceSummary_inst_l_tax_dvalid,
    l_tax_last => PriceSummary_inst_l_tax_last,
    l_tax => PriceSummary_inst_l_tax,
    l_returnflag_valid => PriceSummary_inst_l_returnflag_valid,
    l_returnflag_ready => PriceSummary_inst_l_returnflag_ready,
    l_returnflag_dvalid => PriceSummary_inst_l_returnflag_dvalid,
    l_returnflag_last => PriceSummary_inst_l_returnflag_last,
    l_returnflag_length => PriceSummary_inst_l_returnflag_length,
    l_returnflag_count => PriceSummary_inst_l_returnflag_count,
    l_returnflag_chars_valid => PriceSummary_inst_l_returnflag_chars_valid,
    l_returnflag_chars_ready => PriceSummary_inst_l_returnflag_chars_ready,
    l_returnflag_chars_dvalid => PriceSummary_inst_l_returnflag_chars_dvalid,
    l_returnflag_chars_last => PriceSummary_inst_l_returnflag_chars_last,
    l_returnflag_chars => PriceSummary_inst_l_returnflag_chars,
    l_returnflag_chars_count => PriceSummary_inst_l_returnflag_chars_count,
    l_linestatus_valid => PriceSummary_inst_l_linestatus_valid,
    l_linestatus_ready => PriceSummary_inst_l_linestatus_ready,
    l_linestatus_dvalid => PriceSummary_inst_l_linestatus_dvalid,
    l_linestatus_last => PriceSummary_inst_l_linestatus_last,
    l_linestatus_length => PriceSummary_inst_l_linestatus_length,
    l_linestatus_count => PriceSummary_inst_l_linestatus_count,
    l_linestatus_chars_valid => PriceSummary_inst_l_linestatus_chars_valid,
    l_linestatus_chars_ready => PriceSummary_inst_l_linestatus_chars_ready,
    l_linestatus_chars_dvalid => PriceSummary_inst_l_linestatus_chars_dvalid,
    l_linestatus_chars_last => PriceSummary_inst_l_linestatus_chars_last,
    l_linestatus_chars => PriceSummary_inst_l_linestatus_chars,
    l_linestatus_chars_count => PriceSummary_inst_l_linestatus_chars_count,
    l_shipdate_valid => PriceSummary_inst_l_shipdate_valid,
    l_shipdate_ready => PriceSummary_inst_l_shipdate_ready,
    l_shipdate_dvalid => PriceSummary_inst_l_shipdate_dvalid,
    l_shipdate_last => PriceSummary_inst_l_shipdate_last,
    l_shipdate => PriceSummary_inst_l_shipdate,
    l_quantity_unl_valid => PriceSummary_inst_l_quantity_unl_valid,
    l_quantity_unl_ready => PriceSummary_inst_l_quantity_unl_ready,
    l_quantity_unl_tag => PriceSummary_inst_l_quantity_unl_tag,
    l_extendedprice_unl_valid => PriceSummary_inst_l_extendedprice_unl_valid,
    l_extendedprice_unl_ready => PriceSummary_inst_l_extendedprice_unl_ready,
    l_extendedprice_unl_tag => PriceSummary_inst_l_extendedprice_unl_tag,
    l_discount_unl_valid => PriceSummary_inst_l_discount_unl_valid,
    l_discount_unl_ready => PriceSummary_inst_l_discount_unl_ready,
    l_discount_unl_tag => PriceSummary_inst_l_discount_unl_tag,
    l_tax_unl_valid => PriceSummary_inst_l_tax_unl_valid,
    l_tax_unl_ready => PriceSummary_inst_l_tax_unl_ready,
    l_tax_unl_tag => PriceSummary_inst_l_tax_unl_tag,
    l_returnflag_unl_valid => PriceSummary_inst_l_returnflag_unl_valid,
    l_returnflag_unl_ready => PriceSummary_inst_l_returnflag_unl_ready,
    l_returnflag_unl_tag => PriceSummary_inst_l_returnflag_unl_tag,
    l_linestatus_unl_valid => PriceSummary_inst_l_linestatus_unl_valid,
    l_linestatus_unl_ready => PriceSummary_inst_l_linestatus_unl_ready,
    l_linestatus_unl_tag => PriceSummary_inst_l_linestatus_unl_tag,
    l_shipdate_unl_valid => PriceSummary_inst_l_shipdate_unl_valid,
    l_shipdate_unl_ready => PriceSummary_inst_l_shipdate_unl_ready,
    l_shipdate_unl_tag => PriceSummary_inst_l_shipdate_unl_tag,
    l_quantity_cmd_valid => PriceSummary_inst_l_quantity_cmd_valid,
    l_quantity_cmd_ready => PriceSummary_inst_l_quantity_cmd_ready,
    l_quantity_cmd_firstIdx => PriceSummary_inst_l_quantity_cmd_firstIdx,
    l_quantity_cmd_lastIdx => PriceSummary_inst_l_quantity_cmd_lastIdx,
    l_quantity_cmd_tag => PriceSummary_inst_l_quantity_cmd_tag,
    l_extendedprice_cmd_valid => PriceSummary_inst_l_extendedprice_cmd_valid,
    l_extendedprice_cmd_ready => PriceSummary_inst_l_extendedprice_cmd_ready,
    l_extendedprice_cmd_firstIdx => PriceSummary_inst_l_extendedprice_cmd_firstIdx,
    l_extendedprice_cmd_lastIdx => PriceSummary_inst_l_extendedprice_cmd_lastIdx,
    l_extendedprice_cmd_tag => PriceSummary_inst_l_extendedprice_cmd_tag,
    l_discount_cmd_valid => PriceSummary_inst_l_discount_cmd_valid,
    l_discount_cmd_ready => PriceSummary_inst_l_discount_cmd_ready,
    l_discount_cmd_firstIdx => PriceSummary_inst_l_discount_cmd_firstIdx,
    l_discount_cmd_lastIdx => PriceSummary_inst_l_discount_cmd_lastIdx,
    l_discount_cmd_tag => PriceSummary_inst_l_discount_cmd_tag,
    l_tax_cmd_valid => PriceSummary_inst_l_tax_cmd_valid,
    l_tax_cmd_ready => PriceSummary_inst_l_tax_cmd_ready,
    l_tax_cmd_firstIdx => PriceSummary_inst_l_tax_cmd_firstIdx,
    l_tax_cmd_lastIdx => PriceSummary_inst_l_tax_cmd_lastIdx,
    l_tax_cmd_tag => PriceSummary_inst_l_tax_cmd_tag,
    l_returnflag_cmd_valid => PriceSummary_inst_l_returnflag_cmd_valid,
    l_returnflag_cmd_ready => PriceSummary_inst_l_returnflag_cmd_ready,
    l_returnflag_cmd_firstIdx => PriceSummary_inst_l_returnflag_cmd_firstIdx,
    l_returnflag_cmd_lastIdx => PriceSummary_inst_l_returnflag_cmd_lastIdx,
    l_returnflag_cmd_tag => PriceSummary_inst_l_returnflag_cmd_tag,
    l_linestatus_cmd_valid => PriceSummary_inst_l_linestatus_cmd_valid,
    l_linestatus_cmd_ready => PriceSummary_inst_l_linestatus_cmd_ready,
    l_linestatus_cmd_firstIdx => PriceSummary_inst_l_linestatus_cmd_firstIdx,
    l_linestatus_cmd_lastIdx => PriceSummary_inst_l_linestatus_cmd_lastIdx,
    l_linestatus_cmd_tag => PriceSummary_inst_l_linestatus_cmd_tag,
    l_shipdate_cmd_valid => PriceSummary_inst_l_shipdate_cmd_valid,
    l_shipdate_cmd_ready => PriceSummary_inst_l_shipdate_cmd_ready,
    l_shipdate_cmd_firstIdx => PriceSummary_inst_l_shipdate_cmd_firstIdx,
    l_shipdate_cmd_lastIdx => PriceSummary_inst_l_shipdate_cmd_lastIdx,
    l_shipdate_cmd_tag => PriceSummary_inst_l_shipdate_cmd_tag,
    l_returnflag_o_valid => PriceSummaryWriter_inst_l_returnflag_o_valid,
    l_returnflag_o_ready => PriceSummaryWriter_inst_l_returnflag_o_ready,
    l_returnflag_o_dvalid => PriceSummaryWriter_inst_l_returnflag_o_dvalid,
    l_returnflag_o_last => PriceSummaryWriter_inst_l_returnflag_o_last,
    l_returnflag_o_length => PriceSummaryWriter_inst_l_returnflag_o_length,
    l_returnflag_o_count => PriceSummaryWriter_inst_l_returnflag_o_count,
    l_returnflag_o_chars_valid => PriceSummaryWriter_inst_l_returnflag_o_chars_valid,
    l_returnflag_o_chars_ready => PriceSummaryWriter_inst_l_returnflag_o_chars_ready,
    l_returnflag_o_chars_dvalid => PriceSummaryWriter_inst_l_returnflag_o_chars_dvalid,
    l_returnflag_o_chars_last => PriceSummaryWriter_inst_l_returnflag_o_chars_last,
    l_returnflag_o_chars => PriceSummaryWriter_inst_l_returnflag_o_chars,
    l_returnflag_o_chars_count => PriceSummaryWriter_inst_l_returnflag_o_chars_count,
    l_linestatus_o_valid => PriceSummaryWriter_inst_l_linestatus_o_valid,
    l_linestatus_o_ready => PriceSummaryWriter_inst_l_linestatus_o_ready,
    l_linestatus_o_dvalid => PriceSummaryWriter_inst_l_linestatus_o_dvalid,
    l_linestatus_o_last => PriceSummaryWriter_inst_l_linestatus_o_last,
    l_linestatus_o_length => PriceSummaryWriter_inst_l_linestatus_o_length,
    l_linestatus_o_count => PriceSummaryWriter_inst_l_linestatus_o_count,
    l_linestatus_o_chars_valid => PriceSummaryWriter_inst_l_linestatus_o_chars_valid,
    l_linestatus_o_chars_ready => PriceSummaryWriter_inst_l_linestatus_o_chars_ready,
    l_linestatus_o_chars_dvalid => PriceSummaryWriter_inst_l_linestatus_o_chars_dvalid,
    l_linestatus_o_chars_last => PriceSummaryWriter_inst_l_linestatus_o_chars_last,
    l_linestatus_o_chars => PriceSummaryWriter_inst_l_linestatus_o_chars,
    l_linestatus_o_chars_count => PriceSummaryWriter_inst_l_linestatus_o_chars_count,
    l_sum_qty_valid => PriceSummaryWriter_inst_l_sum_qty_valid,
    l_sum_qty_ready => PriceSummaryWriter_inst_l_sum_qty_ready,
    l_sum_qty_dvalid => PriceSummaryWriter_inst_l_sum_qty_dvalid,
    l_sum_qty_last => PriceSummaryWriter_inst_l_sum_qty_last,
    l_sum_qty => PriceSummaryWriter_inst_l_sum_qty,
    l_sum_base_price_valid => PriceSummaryWriter_inst_l_sum_base_price_valid,
    l_sum_base_price_ready => PriceSummaryWriter_inst_l_sum_base_price_ready,
    l_sum_base_price_dvalid => PriceSummaryWriter_inst_l_sum_base_price_dvalid,
    l_sum_base_price_last => PriceSummaryWriter_inst_l_sum_base_price_last,
    l_sum_base_price => PriceSummaryWriter_inst_l_sum_base_price,
    l_sum_disc_price_valid => PriceSummaryWriter_inst_l_sum_disc_price_valid,
    l_sum_disc_price_ready => PriceSummaryWriter_inst_l_sum_disc_price_ready,
    l_sum_disc_price_dvalid => PriceSummaryWriter_inst_l_sum_disc_price_dvalid,
    l_sum_disc_price_last => PriceSummaryWriter_inst_l_sum_disc_price_last,
    l_sum_disc_price => PriceSummaryWriter_inst_l_sum_disc_price,
    l_sum_charge_valid => PriceSummaryWriter_inst_l_sum_charge_valid,
    l_sum_charge_ready => PriceSummaryWriter_inst_l_sum_charge_ready,
    l_sum_charge_dvalid => PriceSummaryWriter_inst_l_sum_charge_dvalid,
    l_sum_charge_last => PriceSummaryWriter_inst_l_sum_charge_last,
    l_sum_charge => PriceSummaryWriter_inst_l_sum_charge,
    l_avg_qty_valid => PriceSummaryWriter_inst_l_avg_qty_valid,
    l_avg_qty_ready => PriceSummaryWriter_inst_l_avg_qty_ready,
    l_avg_qty_dvalid => PriceSummaryWriter_inst_l_avg_qty_dvalid,
    l_avg_qty_last => PriceSummaryWriter_inst_l_avg_qty_last,
    l_avg_qty => PriceSummaryWriter_inst_l_avg_qty,
    l_avg_price_valid => PriceSummaryWriter_inst_l_avg_price_valid,
    l_avg_price_ready => PriceSummaryWriter_inst_l_avg_price_ready,
    l_avg_price_dvalid => PriceSummaryWriter_inst_l_avg_price_dvalid,
    l_avg_price_last => PriceSummaryWriter_inst_l_avg_price_last,
    l_avg_price => PriceSummaryWriter_inst_l_avg_price,
    l_avg_disc_valid => PriceSummaryWriter_inst_l_avg_disc_valid,
    l_avg_disc_ready => PriceSummaryWriter_inst_l_avg_disc_ready,
    l_avg_disc_dvalid => PriceSummaryWriter_inst_l_avg_disc_dvalid,
    l_avg_disc_last => PriceSummaryWriter_inst_l_avg_disc_last,
    l_avg_disc => PriceSummaryWriter_inst_l_avg_disc,
    l_count_order_valid => PriceSummaryWriter_inst_l_count_order_valid,
    l_count_order_ready => PriceSummaryWriter_inst_l_count_order_ready,
    l_count_order_dvalid => PriceSummaryWriter_inst_l_count_order_dvalid,
    l_count_order_last => PriceSummaryWriter_inst_l_count_order_last,
    l_count_order => PriceSummaryWriter_inst_l_count_order,
    l_returnflag_o_unl_valid => PriceSummaryWriter_inst_l_returnflag_o_unl_valid,
    l_returnflag_o_unl_ready => PriceSummaryWriter_inst_l_returnflag_o_unl_ready,
    l_returnflag_o_unl_tag => PriceSummaryWriter_inst_l_returnflag_o_unl_tag,
    l_linestatus_o_unl_valid => PriceSummaryWriter_inst_l_linestatus_o_unl_valid,
    l_linestatus_o_unl_ready => PriceSummaryWriter_inst_l_linestatus_o_unl_ready,
    l_linestatus_o_unl_tag => PriceSummaryWriter_inst_l_linestatus_o_unl_tag,
    l_sum_qty_unl_valid => PriceSummaryWriter_inst_l_sum_qty_unl_valid,
    l_sum_qty_unl_ready => PriceSummaryWriter_inst_l_sum_qty_unl_ready,
    l_sum_qty_unl_tag => PriceSummaryWriter_inst_l_sum_qty_unl_tag,
    l_sum_base_price_unl_valid => PriceSummaryWriter_inst_l_sum_base_price_unl_valid,
    l_sum_base_price_unl_ready => PriceSummaryWriter_inst_l_sum_base_price_unl_ready,
    l_sum_base_price_unl_tag => PriceSummaryWriter_inst_l_sum_base_price_unl_tag,
    l_sum_disc_price_unl_valid => PriceSummaryWriter_inst_l_sum_disc_price_unl_valid,
    l_sum_disc_price_unl_ready => PriceSummaryWriter_inst_l_sum_disc_price_unl_ready,
    l_sum_disc_price_unl_tag => PriceSummaryWriter_inst_l_sum_disc_price_unl_tag,
    l_sum_charge_unl_valid => PriceSummaryWriter_inst_l_sum_charge_unl_valid,
    l_sum_charge_unl_ready => PriceSummaryWriter_inst_l_sum_charge_unl_ready,
    l_sum_charge_unl_tag => PriceSummaryWriter_inst_l_sum_charge_unl_tag,
    l_avg_qty_unl_valid => PriceSummaryWriter_inst_l_avg_qty_unl_valid,
    l_avg_qty_unl_ready => PriceSummaryWriter_inst_l_avg_qty_unl_ready,
    l_avg_qty_unl_tag => PriceSummaryWriter_inst_l_avg_qty_unl_tag,
    l_avg_price_unl_valid => PriceSummaryWriter_inst_l_avg_price_unl_valid,
    l_avg_price_unl_ready => PriceSummaryWriter_inst_l_avg_price_unl_ready,
    l_avg_price_unl_tag => PriceSummaryWriter_inst_l_avg_price_unl_tag,
    l_avg_disc_unl_valid => PriceSummaryWriter_inst_l_avg_disc_unl_valid,
    l_avg_disc_unl_ready => PriceSummaryWriter_inst_l_avg_disc_unl_ready,
    l_avg_disc_unl_tag => PriceSummaryWriter_inst_l_avg_disc_unl_tag,
    l_count_order_unl_valid => PriceSummaryWriter_inst_l_count_order_unl_valid,
    l_count_order_unl_ready => PriceSummaryWriter_inst_l_count_order_unl_ready,
    l_count_order_unl_tag => PriceSummaryWriter_inst_l_count_order_unl_tag,
    l_returnflag_o_cmd_valid => PriceSummaryWriter_inst_l_returnflag_o_cmd_valid,
    l_returnflag_o_cmd_ready => PriceSummaryWriter_inst_l_returnflag_o_cmd_ready,
    l_returnflag_o_cmd_firstIdx => PriceSummaryWriter_inst_l_returnflag_o_cmd_firstIdx,
    l_returnflag_o_cmd_lastIdx => PriceSummaryWriter_inst_l_returnflag_o_cmd_lastIdx,
    l_returnflag_o_cmd_tag => PriceSummaryWriter_inst_l_returnflag_o_cmd_tag,
    l_linestatus_o_cmd_valid => PriceSummaryWriter_inst_l_linestatus_o_cmd_valid,
    l_linestatus_o_cmd_ready => PriceSummaryWriter_inst_l_linestatus_o_cmd_ready,
    l_linestatus_o_cmd_firstIdx => PriceSummaryWriter_inst_l_linestatus_o_cmd_firstIdx,
    l_linestatus_o_cmd_lastIdx => PriceSummaryWriter_inst_l_linestatus_o_cmd_lastIdx,
    l_linestatus_o_cmd_tag => PriceSummaryWriter_inst_l_linestatus_o_cmd_tag,
    l_sum_qty_cmd_valid => PriceSummaryWriter_inst_l_sum_qty_cmd_valid,
    l_sum_qty_cmd_ready => PriceSummaryWriter_inst_l_sum_qty_cmd_ready,
    l_sum_qty_cmd_firstIdx => PriceSummaryWriter_inst_l_sum_qty_cmd_firstIdx,
    l_sum_qty_cmd_lastIdx => PriceSummaryWriter_inst_l_sum_qty_cmd_lastIdx,
    l_sum_qty_cmd_tag => PriceSummaryWriter_inst_l_sum_qty_cmd_tag,
    l_sum_base_price_cmd_valid => PriceSummaryWriter_inst_l_sum_base_price_cmd_valid,
    l_sum_base_price_cmd_ready => PriceSummaryWriter_inst_l_sum_base_price_cmd_ready,
    l_sum_base_price_cmd_firstIdx => PriceSummaryWriter_inst_l_sum_base_price_cmd_firstIdx,
    l_sum_base_price_cmd_lastIdx => PriceSummaryWriter_inst_l_sum_base_price_cmd_lastIdx,
    l_sum_base_price_cmd_tag => PriceSummaryWriter_inst_l_sum_base_price_cmd_tag,
    l_sum_disc_price_cmd_valid => PriceSummaryWriter_inst_l_sum_disc_price_cmd_valid,
    l_sum_disc_price_cmd_ready => PriceSummaryWriter_inst_l_sum_disc_price_cmd_ready,
    l_sum_disc_price_cmd_firstIdx => PriceSummaryWriter_inst_l_sum_disc_price_cmd_firstIdx,
    l_sum_disc_price_cmd_lastIdx => PriceSummaryWriter_inst_l_sum_disc_price_cmd_lastIdx,
    l_sum_disc_price_cmd_tag => PriceSummaryWriter_inst_l_sum_disc_price_cmd_tag,
    l_sum_charge_cmd_valid => PriceSummaryWriter_inst_l_sum_charge_cmd_valid,
    l_sum_charge_cmd_ready => PriceSummaryWriter_inst_l_sum_charge_cmd_ready,
    l_sum_charge_cmd_firstIdx => PriceSummaryWriter_inst_l_sum_charge_cmd_firstIdx,
    l_sum_charge_cmd_lastIdx => PriceSummaryWriter_inst_l_sum_charge_cmd_lastIdx,
    l_sum_charge_cmd_tag => PriceSummaryWriter_inst_l_sum_charge_cmd_tag,
    l_avg_qty_cmd_valid => PriceSummaryWriter_inst_l_avg_qty_cmd_valid,
    l_avg_qty_cmd_ready => PriceSummaryWriter_inst_l_avg_qty_cmd_ready,
    l_avg_qty_cmd_firstIdx => PriceSummaryWriter_inst_l_avg_qty_cmd_firstIdx,
    l_avg_qty_cmd_lastIdx => PriceSummaryWriter_inst_l_avg_qty_cmd_lastIdx,
    l_avg_qty_cmd_tag => PriceSummaryWriter_inst_l_avg_qty_cmd_tag,
    l_avg_price_cmd_valid => PriceSummaryWriter_inst_l_avg_price_cmd_valid,
    l_avg_price_cmd_ready => PriceSummaryWriter_inst_l_avg_price_cmd_ready,
    l_avg_price_cmd_firstIdx => PriceSummaryWriter_inst_l_avg_price_cmd_firstIdx,
    l_avg_price_cmd_lastIdx => PriceSummaryWriter_inst_l_avg_price_cmd_lastIdx,
    l_avg_price_cmd_tag => PriceSummaryWriter_inst_l_avg_price_cmd_tag,
    l_avg_disc_cmd_valid => PriceSummaryWriter_inst_l_avg_disc_cmd_valid,
    l_avg_disc_cmd_ready => PriceSummaryWriter_inst_l_avg_disc_cmd_ready,
    l_avg_disc_cmd_firstIdx => PriceSummaryWriter_inst_l_avg_disc_cmd_firstIdx,
    l_avg_disc_cmd_lastIdx => PriceSummaryWriter_inst_l_avg_disc_cmd_lastIdx,
    l_avg_disc_cmd_tag => PriceSummaryWriter_inst_l_avg_disc_cmd_tag,
    l_count_order_cmd_valid => PriceSummaryWriter_inst_l_count_order_cmd_valid,
    l_count_order_cmd_ready => PriceSummaryWriter_inst_l_count_order_cmd_ready,
    l_count_order_cmd_firstIdx => PriceSummaryWriter_inst_l_count_order_cmd_firstIdx,
    l_count_order_cmd_lastIdx => PriceSummaryWriter_inst_l_count_order_cmd_lastIdx,
    l_count_order_cmd_tag => PriceSummaryWriter_inst_l_count_order_cmd_tag,
    start => PriceSummary_inst_start,
    stop => PriceSummary_inst_stop,
    reset => PriceSummary_inst_reset,
    idle => PriceSummary_inst_idle,
    busy => PriceSummary_inst_busy,
    done => PriceSummary_inst_done,
    result => PriceSummary_inst_result,
    l_firstidx => PriceSummary_inst_l_firstidx,
    l_lastidx => PriceSummary_inst_l_lastidx,
    rhigh => PriceSummary_inst_rhigh,
    rlow => PriceSummary_inst_rlow,
    status_1 => PriceSummary_inst_status_1,
    status_2 => PriceSummary_inst_status_2,
    r1 => PriceSummary_inst_r1,
    r2 => PriceSummary_inst_r2,
    r3 => PriceSummary_inst_r3,
    r4 => PriceSummary_inst_r4,
    r5 => PriceSummary_inst_r5,
    r6 => PriceSummary_inst_r6,
    r7 => PriceSummary_inst_r7,
    r8 => PriceSummary_inst_r8
  );

  mmio_inst : mmio
  PORT MAP(
    kcd_clk => kcd_clk,
    kcd_reset => kcd_reset,
    f_start_data => mmio_inst_f_start_data,
    f_stop_data => mmio_inst_f_stop_data,
    f_reset_data => mmio_inst_f_reset_data,
    f_idle_write_data => mmio_inst_f_idle_write_data,
    f_busy_write_data => mmio_inst_f_busy_write_data,
    f_done_write_data => mmio_inst_f_done_write_data,
    f_result_write_data => mmio_inst_f_result_write_data,
    f_l_firstidx_data => mmio_inst_f_l_firstidx_data,
    f_l_lastidx_data => mmio_inst_f_l_lastidx_data,
    f_l_quantity_values_data => mmio_inst_f_l_quantity_values_data,
    f_l_extendedprice_values_data => mmio_inst_f_l_extendedprice_values_data,
    f_l_discount_values_data => mmio_inst_f_l_discount_values_data,
    f_l_tax_values_data => mmio_inst_f_l_tax_values_data,
    f_l_returnflag_offsets_data => mmio_inst_f_l_returnflag_offsets_data,
    f_l_returnflag_values_data => mmio_inst_f_l_returnflag_values_data,
    f_l_linestatus_offsets_data => mmio_inst_f_l_linestatus_offsets_data,
    f_l_linestatus_values_data => mmio_inst_f_l_linestatus_values_data,
    f_l_shipdate_values_data => mmio_inst_f_l_shipdate_values_data,
    l_returnflag_o_valid => PriceSummaryWriter_inst_l_returnflag_o_valid,
    l_returnflag_o_ready => PriceSummaryWriter_inst_l_returnflag_o_ready,
    l_returnflag_o_dvalid => PriceSummaryWriter_inst_l_returnflag_o_dvalid,
    l_returnflag_o_last => PriceSummaryWriter_inst_l_returnflag_o_last,
    l_returnflag_o_length => PriceSummaryWriter_inst_l_returnflag_o_length,
    l_returnflag_o_count => PriceSummaryWriter_inst_l_returnflag_o_count,
    l_returnflag_o_chars_valid => PriceSummaryWriter_inst_l_returnflag_o_chars_valid,
    l_returnflag_o_chars_ready => PriceSummaryWriter_inst_l_returnflag_o_chars_ready,
    l_returnflag_o_chars_dvalid => PriceSummaryWriter_inst_l_returnflag_o_chars_dvalid,
    l_returnflag_o_chars_last => PriceSummaryWriter_inst_l_returnflag_o_chars_last,
    l_returnflag_o_chars => PriceSummaryWriter_inst_l_returnflag_o_chars,
    l_returnflag_o_chars_count => PriceSummaryWriter_inst_l_returnflag_o_chars_count,
    l_linestatus_o_valid => PriceSummaryWriter_inst_l_linestatus_o_valid,
    l_linestatus_o_ready => PriceSummaryWriter_inst_l_linestatus_o_ready,
    l_linestatus_o_dvalid => PriceSummaryWriter_inst_l_linestatus_o_dvalid,
    l_linestatus_o_last => PriceSummaryWriter_inst_l_linestatus_o_last,
    l_linestatus_o_length => PriceSummaryWriter_inst_l_linestatus_o_length,
    l_linestatus_o_count => PriceSummaryWriter_inst_l_linestatus_o_count,
    l_linestatus_o_chars_valid => PriceSummaryWriter_inst_l_linestatus_o_chars_valid,
    l_linestatus_o_chars_ready => PriceSummaryWriter_inst_l_linestatus_o_chars_ready,
    l_linestatus_o_chars_dvalid => PriceSummaryWriter_inst_l_linestatus_o_chars_dvalid,
    l_linestatus_o_chars_last => PriceSummaryWriter_inst_l_linestatus_o_chars_last,
    l_linestatus_o_chars => PriceSummaryWriter_inst_l_linestatus_o_chars,
    l_linestatus_o_chars_count => PriceSummaryWriter_inst_l_linestatus_o_chars_count,
    l_sum_qty_valid => PriceSummaryWriter_inst_l_sum_qty_valid,
    l_sum_qty_ready => PriceSummaryWriter_inst_l_sum_qty_ready,
    l_sum_qty_dvalid => PriceSummaryWriter_inst_l_sum_qty_dvalid,
    l_sum_qty_last => PriceSummaryWriter_inst_l_sum_qty_last,
    l_sum_qty => PriceSummaryWriter_inst_l_sum_qty,
    l_sum_base_price_valid => PriceSummaryWriter_inst_l_sum_base_price_valid,
    l_sum_base_price_ready => PriceSummaryWriter_inst_l_sum_base_price_ready,
    l_sum_base_price_dvalid => PriceSummaryWriter_inst_l_sum_base_price_dvalid,
    l_sum_base_price_last => PriceSummaryWriter_inst_l_sum_base_price_last,
    l_sum_base_price => PriceSummaryWriter_inst_l_sum_base_price,
    l_sum_disc_price_valid => PriceSummaryWriter_inst_l_sum_disc_price_valid,
    l_sum_disc_price_ready => PriceSummaryWriter_inst_l_sum_disc_price_ready,
    l_sum_disc_price_dvalid => PriceSummaryWriter_inst_l_sum_disc_price_dvalid,
    l_sum_disc_price_last => PriceSummaryWriter_inst_l_sum_disc_price_last,
    l_sum_disc_price => PriceSummaryWriter_inst_l_sum_disc_price,
    l_sum_charge_valid => PriceSummaryWriter_inst_l_sum_charge_valid,
    l_sum_charge_ready => PriceSummaryWriter_inst_l_sum_charge_ready,
    l_sum_charge_dvalid => PriceSummaryWriter_inst_l_sum_charge_dvalid,
    l_sum_charge_last => PriceSummaryWriter_inst_l_sum_charge_last,
    l_sum_charge => PriceSummaryWriter_inst_l_sum_charge,
    l_avg_qty_valid => PriceSummaryWriter_inst_l_avg_qty_valid,
    l_avg_qty_ready => PriceSummaryWriter_inst_l_avg_qty_ready,
    l_avg_qty_dvalid => PriceSummaryWriter_inst_l_avg_qty_dvalid,
    l_avg_qty_last => PriceSummaryWriter_inst_l_avg_qty_last,
    l_avg_qty => PriceSummaryWriter_inst_l_avg_qty,
    l_avg_price_valid => PriceSummaryWriter_inst_l_avg_price_valid,
    l_avg_price_ready => PriceSummaryWriter_inst_l_avg_price_ready,
    l_avg_price_dvalid => PriceSummaryWriter_inst_l_avg_price_dvalid,
    l_avg_price_last => PriceSummaryWriter_inst_l_avg_price_last,
    l_avg_price => PriceSummaryWriter_inst_l_avg_price,
    l_avg_disc_valid => PriceSummaryWriter_inst_l_avg_disc_valid,
    l_avg_disc_ready => PriceSummaryWriter_inst_l_avg_disc_ready,
    l_avg_disc_dvalid => PriceSummaryWriter_inst_l_avg_disc_dvalid,
    l_avg_disc_last => PriceSummaryWriter_inst_l_avg_disc_last,
    l_avg_disc => PriceSummaryWriter_inst_l_avg_disc,
    l_count_order_valid => PriceSummaryWriter_inst_l_count_order_valid,
    l_count_order_ready => PriceSummaryWriter_inst_l_count_order_ready,
    l_count_order_dvalid => PriceSummaryWriter_inst_l_count_order_dvalid,
    l_count_order_last => PriceSummaryWriter_inst_l_count_order_last,
    l_count_order => PriceSummaryWriter_inst_l_count_order,
    l_returnflag_o_unl_valid => PriceSummaryWriter_inst_l_returnflag_o_unl_valid,
    l_returnflag_o_unl_ready => PriceSummaryWriter_inst_l_returnflag_o_unl_ready,
    l_returnflag_o_unl_tag => PriceSummaryWriter_inst_l_returnflag_o_unl_tag,
    l_linestatus_o_unl_valid => PriceSummaryWriter_inst_l_linestatus_o_unl_valid,
    l_linestatus_o_unl_ready => PriceSummaryWriter_inst_l_linestatus_o_unl_ready,
    l_linestatus_o_unl_tag => PriceSummaryWriter_inst_l_linestatus_o_unl_tag,
    l_sum_qty_unl_valid => PriceSummaryWriter_inst_l_sum_qty_unl_valid,
    l_sum_qty_unl_ready => PriceSummaryWriter_inst_l_sum_qty_unl_ready,
    l_sum_qty_unl_tag => PriceSummaryWriter_inst_l_sum_qty_unl_tag,
    l_sum_base_price_unl_valid => PriceSummaryWriter_inst_l_sum_base_price_unl_valid,
    l_sum_base_price_unl_ready => PriceSummaryWriter_inst_l_sum_base_price_unl_ready,
    l_sum_base_price_unl_tag => PriceSummaryWriter_inst_l_sum_base_price_unl_tag,
    l_sum_disc_price_unl_valid => PriceSummaryWriter_inst_l_sum_disc_price_unl_valid,
    l_sum_disc_price_unl_ready => PriceSummaryWriter_inst_l_sum_disc_price_unl_ready,
    l_sum_disc_price_unl_tag => PriceSummaryWriter_inst_l_sum_disc_price_unl_tag,
    l_sum_charge_unl_valid => PriceSummaryWriter_inst_l_sum_charge_unl_valid,
    l_sum_charge_unl_ready => PriceSummaryWriter_inst_l_sum_charge_unl_ready,
    l_sum_charge_unl_tag => PriceSummaryWriter_inst_l_sum_charge_unl_tag,
    l_avg_qty_unl_valid => PriceSummaryWriter_inst_l_avg_qty_unl_valid,
    l_avg_qty_unl_ready => PriceSummaryWriter_inst_l_avg_qty_unl_ready,
    l_avg_qty_unl_tag => PriceSummaryWriter_inst_l_avg_qty_unl_tag,
    l_avg_price_unl_valid => PriceSummaryWriter_inst_l_avg_price_unl_valid,
    l_avg_price_unl_ready => PriceSummaryWriter_inst_l_avg_price_unl_ready,
    l_avg_price_unl_tag => PriceSummaryWriter_inst_l_avg_price_unl_tag,
    l_avg_disc_unl_valid => PriceSummaryWriter_inst_l_avg_disc_unl_valid,
    l_avg_disc_unl_ready => PriceSummaryWriter_inst_l_avg_disc_unl_ready,
    l_avg_disc_unl_tag => PriceSummaryWriter_inst_l_avg_disc_unl_tag,
    l_count_order_unl_valid => PriceSummaryWriter_inst_l_count_order_unl_valid,
    l_count_order_unl_ready => PriceSummaryWriter_inst_l_count_order_unl_ready,
    l_count_order_unl_tag => PriceSummaryWriter_inst_l_count_order_unl_tag,
    l_returnflag_o_cmd_valid => PriceSummaryWriter_inst_l_returnflag_o_cmd_valid,
    l_returnflag_o_cmd_ready => PriceSummaryWriter_inst_l_returnflag_o_cmd_ready,
    l_returnflag_o_cmd_firstIdx => PriceSummaryWriter_inst_l_returnflag_o_cmd_firstIdx,
    l_returnflag_o_cmd_lastIdx => PriceSummaryWriter_inst_l_returnflag_o_cmd_lastIdx,
    l_returnflag_o_cmd_tag => PriceSummaryWriter_inst_l_returnflag_o_cmd_tag,
    l_linestatus_o_cmd_valid => PriceSummaryWriter_inst_l_linestatus_o_cmd_valid,
    l_linestatus_o_cmd_ready => PriceSummaryWriter_inst_l_linestatus_o_cmd_ready,
    l_linestatus_o_cmd_firstIdx => PriceSummaryWriter_inst_l_linestatus_o_cmd_firstIdx,
    l_linestatus_o_cmd_lastIdx => PriceSummaryWriter_inst_l_linestatus_o_cmd_lastIdx,
    l_linestatus_o_cmd_tag => PriceSummaryWriter_inst_l_linestatus_o_cmd_tag,
    l_sum_qty_cmd_valid => PriceSummaryWriter_inst_l_sum_qty_cmd_valid,
    l_sum_qty_cmd_ready => PriceSummaryWriter_inst_l_sum_qty_cmd_ready,
    l_sum_qty_cmd_firstIdx => PriceSummaryWriter_inst_l_sum_qty_cmd_firstIdx,
    l_sum_qty_cmd_lastIdx => PriceSummaryWriter_inst_l_sum_qty_cmd_lastIdx,
    l_sum_qty_cmd_tag => PriceSummaryWriter_inst_l_sum_qty_cmd_tag,
    l_sum_base_price_cmd_valid => PriceSummaryWriter_inst_l_sum_base_price_cmd_valid,
    l_sum_base_price_cmd_ready => PriceSummaryWriter_inst_l_sum_base_price_cmd_ready,
    l_sum_base_price_cmd_firstIdx => PriceSummaryWriter_inst_l_sum_base_price_cmd_firstIdx,
    l_sum_base_price_cmd_lastIdx => PriceSummaryWriter_inst_l_sum_base_price_cmd_lastIdx,
    l_sum_base_price_cmd_tag => PriceSummaryWriter_inst_l_sum_base_price_cmd_tag,
    l_sum_disc_price_cmd_valid => PriceSummaryWriter_inst_l_sum_disc_price_cmd_valid,
    l_sum_disc_price_cmd_ready => PriceSummaryWriter_inst_l_sum_disc_price_cmd_ready,
    l_sum_disc_price_cmd_firstIdx => PriceSummaryWriter_inst_l_sum_disc_price_cmd_firstIdx,
    l_sum_disc_price_cmd_lastIdx => PriceSummaryWriter_inst_l_sum_disc_price_cmd_lastIdx,
    l_sum_disc_price_cmd_tag => PriceSummaryWriter_inst_l_sum_disc_price_cmd_tag,
    l_sum_charge_cmd_valid => PriceSummaryWriter_inst_l_sum_charge_cmd_valid,
    l_sum_charge_cmd_ready => PriceSummaryWriter_inst_l_sum_charge_cmd_ready,
    l_sum_charge_cmd_firstIdx => PriceSummaryWriter_inst_l_sum_charge_cmd_firstIdx,
    l_sum_charge_cmd_lastIdx => PriceSummaryWriter_inst_l_sum_charge_cmd_lastIdx,
    l_sum_charge_cmd_tag => PriceSummaryWriter_inst_l_sum_charge_cmd_tag,
    l_avg_qty_cmd_valid => PriceSummaryWriter_inst_l_avg_qty_cmd_valid,
    l_avg_qty_cmd_ready => PriceSummaryWriter_inst_l_avg_qty_cmd_ready,
    l_avg_qty_cmd_firstIdx => PriceSummaryWriter_inst_l_avg_qty_cmd_firstIdx,
    l_avg_qty_cmd_lastIdx => PriceSummaryWriter_inst_l_avg_qty_cmd_lastIdx,
    l_avg_qty_cmd_tag => PriceSummaryWriter_inst_l_avg_qty_cmd_tag,
    l_avg_price_cmd_valid => PriceSummaryWriter_inst_l_avg_price_cmd_valid,
    l_avg_price_cmd_ready => PriceSummaryWriter_inst_l_avg_price_cmd_ready,
    l_avg_price_cmd_firstIdx => PriceSummaryWriter_inst_l_avg_price_cmd_firstIdx,
    l_avg_price_cmd_lastIdx => PriceSummaryWriter_inst_l_avg_price_cmd_lastIdx,
    l_avg_price_cmd_tag => PriceSummaryWriter_inst_l_avg_price_cmd_tag,
    l_avg_disc_cmd_valid => PriceSummaryWriter_inst_l_avg_disc_cmd_valid,
    l_avg_disc_cmd_ready => PriceSummaryWriter_inst_l_avg_disc_cmd_ready,
    l_avg_disc_cmd_firstIdx => PriceSummaryWriter_inst_l_avg_disc_cmd_firstIdx,
    l_avg_disc_cmd_lastIdx => PriceSummaryWriter_inst_l_avg_disc_cmd_lastIdx,
    l_avg_disc_cmd_tag => PriceSummaryWriter_inst_l_avg_disc_cmd_tag,
    l_count_order_cmd_valid => PriceSummaryWriter_inst_l_count_order_cmd_valid,
    l_count_order_cmd_ready => PriceSummaryWriter_inst_l_count_order_cmd_ready,
    l_count_order_cmd_firstIdx => PriceSummaryWriter_inst_l_count_order_cmd_firstIdx,
    l_count_order_cmd_lastIdx => PriceSummaryWriter_inst_l_count_order_cmd_lastIdx,
    l_count_order_cmd_tag => PriceSummaryWriter_inst_l_count_order_cmd_tag,
    f_rhigh_write_data => mmio_inst_f_rhigh_write_data,
    f_rlow_write_data => mmio_inst_f_rlow_write_data,
    f_status_1_write_data => mmio_inst_f_status_1_write_data,
    f_status_2_write_data => mmio_inst_f_status_2_write_data,
    f_r1_write_data => mmio_inst_f_r1_write_data,
    f_r2_write_data => mmio_inst_f_r2_write_data,
    f_r3_write_data => mmio_inst_f_r3_write_data,
    f_r4_write_data => mmio_inst_f_r4_write_data,
    f_r5_write_data => mmio_inst_f_r5_write_data,
    f_r6_write_data => mmio_inst_f_r6_write_data,
    f_r7_write_data => mmio_inst_f_r7_write_data,
    f_r8_write_data => mmio_inst_f_r8_write_data,
    mmio_awvalid => mmio_inst_mmio_awvalid,
    mmio_awready => mmio_inst_mmio_awready,
    mmio_awaddr => mmio_inst_mmio_awaddr,
    mmio_wvalid => mmio_inst_mmio_wvalid,
    mmio_wready => mmio_inst_mmio_wready,
    mmio_wdata => mmio_inst_mmio_wdata,
    mmio_wstrb => mmio_inst_mmio_wstrb,
    mmio_bvalid => mmio_inst_mmio_bvalid,
    mmio_bready => mmio_inst_mmio_bready,
    mmio_bresp => mmio_inst_mmio_bresp,
    mmio_arvalid => mmio_inst_mmio_arvalid,
    mmio_arready => mmio_inst_mmio_arready,
    mmio_araddr => mmio_inst_mmio_araddr,
    mmio_rvalid => mmio_inst_mmio_rvalid,
    mmio_rready => mmio_inst_mmio_rready,
    mmio_rdata => mmio_inst_mmio_rdata,
    mmio_rresp => mmio_inst_mmio_rresp
  );

  l_quantity_cmd_accm_inst : ArrayCmdCtrlMerger
  GENERIC MAP(
    NUM_ADDR => 1,
    BUS_ADDR_WIDTH => L_QUANTITY_BUS_ADDR_WIDTH,
    INDEX_WIDTH => INDEX_WIDTH,
    TAG_WIDTH => TAG_WIDTH
  )
  PORT MAP(
    kernel_cmd_valid => l_quantity_cmd_accm_inst_kernel_cmd_valid,
    kernel_cmd_ready => l_quantity_cmd_accm_inst_kernel_cmd_ready,
    kernel_cmd_firstIdx => l_quantity_cmd_accm_inst_kernel_cmd_firstIdx,
    kernel_cmd_lastIdx => l_quantity_cmd_accm_inst_kernel_cmd_lastIdx,
    kernel_cmd_tag => l_quantity_cmd_accm_inst_kernel_cmd_tag,
    nucleus_cmd_valid => l_quantity_cmd_accm_inst_nucleus_cmd_valid,
    nucleus_cmd_ready => l_quantity_cmd_accm_inst_nucleus_cmd_ready,
    nucleus_cmd_firstIdx => l_quantity_cmd_accm_inst_nucleus_cmd_firstIdx,
    nucleus_cmd_lastIdx => l_quantity_cmd_accm_inst_nucleus_cmd_lastIdx,
    nucleus_cmd_ctrl => l_quantity_cmd_accm_inst_nucleus_cmd_ctrl,
    nucleus_cmd_tag => l_quantity_cmd_accm_inst_nucleus_cmd_tag,
    ctrl => l_quantity_cmd_accm_inst_ctrl
  );

  l_extendedprice_cmd_accm_inst : ArrayCmdCtrlMerger
  GENERIC MAP(
    NUM_ADDR => 1,
    BUS_ADDR_WIDTH => L_EXTENDEDPRICE_BUS_ADDR_WIDTH,
    INDEX_WIDTH => INDEX_WIDTH,
    TAG_WIDTH => TAG_WIDTH
  )
  PORT MAP(
    kernel_cmd_valid => l_extendedprice_cmd_accm_inst_kernel_cmd_valid,
    kernel_cmd_ready => l_extendedprice_cmd_accm_inst_kernel_cmd_ready,
    kernel_cmd_firstIdx => l_extendedprice_cmd_accm_inst_kernel_cmd_firstIdx,
    kernel_cmd_lastIdx => l_extendedprice_cmd_accm_inst_kernel_cmd_lastIdx,
    kernel_cmd_tag => l_extendedprice_cmd_accm_inst_kernel_cmd_tag,
    nucleus_cmd_valid => l_extendedprice_cmd_accm_inst_nucleus_cmd_valid,
    nucleus_cmd_ready => l_extendedprice_cmd_accm_inst_nucleus_cmd_ready,
    nucleus_cmd_firstIdx => l_extendedprice_cmd_accm_inst_nucleus_cmd_firstIdx,
    nucleus_cmd_lastIdx => l_extendedprice_cmd_accm_inst_nucleus_cmd_lastIdx,
    nucleus_cmd_ctrl => l_extendedprice_cmd_accm_inst_nucleus_cmd_ctrl,
    nucleus_cmd_tag => l_extendedprice_cmd_accm_inst_nucleus_cmd_tag,
    ctrl => l_extendedprice_cmd_accm_inst_ctrl
  );

  l_discount_cmd_accm_inst : ArrayCmdCtrlMerger
  GENERIC MAP(
    NUM_ADDR => 1,
    BUS_ADDR_WIDTH => L_DISCOUNT_BUS_ADDR_WIDTH,
    INDEX_WIDTH => INDEX_WIDTH,
    TAG_WIDTH => TAG_WIDTH
  )
  PORT MAP(
    kernel_cmd_valid => l_discount_cmd_accm_inst_kernel_cmd_valid,
    kernel_cmd_ready => l_discount_cmd_accm_inst_kernel_cmd_ready,
    kernel_cmd_firstIdx => l_discount_cmd_accm_inst_kernel_cmd_firstIdx,
    kernel_cmd_lastIdx => l_discount_cmd_accm_inst_kernel_cmd_lastIdx,
    kernel_cmd_tag => l_discount_cmd_accm_inst_kernel_cmd_tag,
    nucleus_cmd_valid => l_discount_cmd_accm_inst_nucleus_cmd_valid,
    nucleus_cmd_ready => l_discount_cmd_accm_inst_nucleus_cmd_ready,
    nucleus_cmd_firstIdx => l_discount_cmd_accm_inst_nucleus_cmd_firstIdx,
    nucleus_cmd_lastIdx => l_discount_cmd_accm_inst_nucleus_cmd_lastIdx,
    nucleus_cmd_ctrl => l_discount_cmd_accm_inst_nucleus_cmd_ctrl,
    nucleus_cmd_tag => l_discount_cmd_accm_inst_nucleus_cmd_tag,
    ctrl => l_discount_cmd_accm_inst_ctrl
  );

  l_tax_cmd_accm_inst : ArrayCmdCtrlMerger
  GENERIC MAP(
    NUM_ADDR => 1,
    BUS_ADDR_WIDTH => L_TAX_BUS_ADDR_WIDTH,
    INDEX_WIDTH => INDEX_WIDTH,
    TAG_WIDTH => TAG_WIDTH
  )
  PORT MAP(
    kernel_cmd_valid => l_tax_cmd_accm_inst_kernel_cmd_valid,
    kernel_cmd_ready => l_tax_cmd_accm_inst_kernel_cmd_ready,
    kernel_cmd_firstIdx => l_tax_cmd_accm_inst_kernel_cmd_firstIdx,
    kernel_cmd_lastIdx => l_tax_cmd_accm_inst_kernel_cmd_lastIdx,
    kernel_cmd_tag => l_tax_cmd_accm_inst_kernel_cmd_tag,
    nucleus_cmd_valid => l_tax_cmd_accm_inst_nucleus_cmd_valid,
    nucleus_cmd_ready => l_tax_cmd_accm_inst_nucleus_cmd_ready,
    nucleus_cmd_firstIdx => l_tax_cmd_accm_inst_nucleus_cmd_firstIdx,
    nucleus_cmd_lastIdx => l_tax_cmd_accm_inst_nucleus_cmd_lastIdx,
    nucleus_cmd_ctrl => l_tax_cmd_accm_inst_nucleus_cmd_ctrl,
    nucleus_cmd_tag => l_tax_cmd_accm_inst_nucleus_cmd_tag,
    ctrl => l_tax_cmd_accm_inst_ctrl
  );

  l_returnflag_cmd_accm_inst : ArrayCmdCtrlMerger
  GENERIC MAP(
    NUM_ADDR => 2,
    BUS_ADDR_WIDTH => L_RETURNFLAG_BUS_ADDR_WIDTH,
    INDEX_WIDTH => INDEX_WIDTH,
    TAG_WIDTH => TAG_WIDTH
  )
  PORT MAP(
    kernel_cmd_valid => l_returnflag_cmd_accm_inst_kernel_cmd_valid,
    kernel_cmd_ready => l_returnflag_cmd_accm_inst_kernel_cmd_ready,
    kernel_cmd_firstIdx => l_returnflag_cmd_accm_inst_kernel_cmd_firstIdx,
    kernel_cmd_lastIdx => l_returnflag_cmd_accm_inst_kernel_cmd_lastIdx,
    kernel_cmd_tag => l_returnflag_cmd_accm_inst_kernel_cmd_tag,
    nucleus_cmd_valid => l_returnflag_cmd_accm_inst_nucleus_cmd_valid,
    nucleus_cmd_ready => l_returnflag_cmd_accm_inst_nucleus_cmd_ready,
    nucleus_cmd_firstIdx => l_returnflag_cmd_accm_inst_nucleus_cmd_firstIdx,
    nucleus_cmd_lastIdx => l_returnflag_cmd_accm_inst_nucleus_cmd_lastIdx,
    nucleus_cmd_ctrl => l_returnflag_cmd_accm_inst_nucleus_cmd_ctrl,
    nucleus_cmd_tag => l_returnflag_cmd_accm_inst_nucleus_cmd_tag,
    ctrl => l_returnflag_cmd_accm_inst_ctrl
  );

  l_linestatus_cmd_accm_inst : ArrayCmdCtrlMerger
  GENERIC MAP(
    NUM_ADDR => 2,
    BUS_ADDR_WIDTH => L_LINESTATUS_BUS_ADDR_WIDTH,
    INDEX_WIDTH => INDEX_WIDTH,
    TAG_WIDTH => TAG_WIDTH
  )
  PORT MAP(
    kernel_cmd_valid => l_linestatus_cmd_accm_inst_kernel_cmd_valid,
    kernel_cmd_ready => l_linestatus_cmd_accm_inst_kernel_cmd_ready,
    kernel_cmd_firstIdx => l_linestatus_cmd_accm_inst_kernel_cmd_firstIdx,
    kernel_cmd_lastIdx => l_linestatus_cmd_accm_inst_kernel_cmd_lastIdx,
    kernel_cmd_tag => l_linestatus_cmd_accm_inst_kernel_cmd_tag,
    nucleus_cmd_valid => l_linestatus_cmd_accm_inst_nucleus_cmd_valid,
    nucleus_cmd_ready => l_linestatus_cmd_accm_inst_nucleus_cmd_ready,
    nucleus_cmd_firstIdx => l_linestatus_cmd_accm_inst_nucleus_cmd_firstIdx,
    nucleus_cmd_lastIdx => l_linestatus_cmd_accm_inst_nucleus_cmd_lastIdx,
    nucleus_cmd_ctrl => l_linestatus_cmd_accm_inst_nucleus_cmd_ctrl,
    nucleus_cmd_tag => l_linestatus_cmd_accm_inst_nucleus_cmd_tag,
    ctrl => l_linestatus_cmd_accm_inst_ctrl
  );

  l_shipdate_cmd_accm_inst : ArrayCmdCtrlMerger
  GENERIC MAP(
    NUM_ADDR => 1,
    BUS_ADDR_WIDTH => L_SHIPDATE_BUS_ADDR_WIDTH,
    INDEX_WIDTH => INDEX_WIDTH,
    TAG_WIDTH => TAG_WIDTH
  )
  PORT MAP(
    kernel_cmd_valid => l_shipdate_cmd_accm_inst_kernel_cmd_valid,
    kernel_cmd_ready => l_shipdate_cmd_accm_inst_kernel_cmd_ready,
    kernel_cmd_firstIdx => l_shipdate_cmd_accm_inst_kernel_cmd_firstIdx,
    kernel_cmd_lastIdx => l_shipdate_cmd_accm_inst_kernel_cmd_lastIdx,
    kernel_cmd_tag => l_shipdate_cmd_accm_inst_kernel_cmd_tag,
    nucleus_cmd_valid => l_shipdate_cmd_accm_inst_nucleus_cmd_valid,
    nucleus_cmd_ready => l_shipdate_cmd_accm_inst_nucleus_cmd_ready,
    nucleus_cmd_firstIdx => l_shipdate_cmd_accm_inst_nucleus_cmd_firstIdx,
    nucleus_cmd_lastIdx => l_shipdate_cmd_accm_inst_nucleus_cmd_lastIdx,
    nucleus_cmd_ctrl => l_shipdate_cmd_accm_inst_nucleus_cmd_ctrl,
    nucleus_cmd_tag => l_shipdate_cmd_accm_inst_nucleus_cmd_tag,
    ctrl => l_shipdate_cmd_accm_inst_ctrl
  );

  l_returnflag_o_cmd_accm_inst : ArrayCmdCtrlMerger
  GENERIC MAP(
    NUM_ADDR => 2,
    BUS_ADDR_WIDTH => L_RETURNFLAG_O_BUS_ADDR_WIDTH,
    INDEX_WIDTH => INDEX_WIDTH,
    TAG_WIDTH => TAG_WIDTH
  )
  PORT MAP(
    kernel_cmd_valid => l_returnflag_o_cmd_accm_inst_kernel_cmd_valid,
    kernel_cmd_ready => l_returnflag_o_cmd_accm_inst_kernel_cmd_ready,
    kernel_cmd_firstIdx => l_returnflag_o_cmd_accm_inst_kernel_cmd_firstIdx,
    kernel_cmd_lastIdx => l_returnflag_o_cmd_accm_inst_kernel_cmd_lastIdx,
    kernel_cmd_tag => l_returnflag_o_cmd_accm_inst_kernel_cmd_tag,
    nucleus_cmd_valid => l_returnflag_o_cmd_accm_inst_nucleus_cmd_valid,
    nucleus_cmd_ready => l_returnflag_o_cmd_accm_inst_nucleus_cmd_ready,
    nucleus_cmd_firstIdx => l_returnflag_o_cmd_accm_inst_nucleus_cmd_firstIdx,
    nucleus_cmd_lastIdx => l_returnflag_o_cmd_accm_inst_nucleus_cmd_lastIdx,
    nucleus_cmd_ctrl => l_returnflag_o_cmd_accm_inst_nucleus_cmd_ctrl,
    nucleus_cmd_tag => l_returnflag_o_cmd_accm_inst_nucleus_cmd_tag,
    ctrl => l_returnflag_o_cmd_accm_inst_ctrl
  );

  l_linestatus_o_cmd_accm_inst : ArrayCmdCtrlMerger
  GENERIC MAP(
    NUM_ADDR => 2,
    BUS_ADDR_WIDTH => L_LINESTATUS_O_BUS_ADDR_WIDTH,
    INDEX_WIDTH => INDEX_WIDTH,
    TAG_WIDTH => TAG_WIDTH
  )
  PORT MAP(
    kernel_cmd_valid => l_linestatus_o_cmd_accm_inst_kernel_cmd_valid,
    kernel_cmd_ready => l_linestatus_o_cmd_accm_inst_kernel_cmd_ready,
    kernel_cmd_firstIdx => l_linestatus_o_cmd_accm_inst_kernel_cmd_firstIdx,
    kernel_cmd_lastIdx => l_linestatus_o_cmd_accm_inst_kernel_cmd_lastIdx,
    kernel_cmd_tag => l_linestatus_o_cmd_accm_inst_kernel_cmd_tag,
    nucleus_cmd_valid => l_linestatus_o_cmd_accm_inst_nucleus_cmd_valid,
    nucleus_cmd_ready => l_linestatus_o_cmd_accm_inst_nucleus_cmd_ready,
    nucleus_cmd_firstIdx => l_linestatus_o_cmd_accm_inst_nucleus_cmd_firstIdx,
    nucleus_cmd_lastIdx => l_linestatus_o_cmd_accm_inst_nucleus_cmd_lastIdx,
    nucleus_cmd_ctrl => l_linestatus_o_cmd_accm_inst_nucleus_cmd_ctrl,
    nucleus_cmd_tag => l_linestatus_o_cmd_accm_inst_nucleus_cmd_tag,
    ctrl => l_linestatus_o_cmd_accm_inst_ctrl
  );

  l_sum_qty_cmd_accm_inst : ArrayCmdCtrlMerger
  GENERIC MAP(
    NUM_ADDR => 1,
    BUS_ADDR_WIDTH => L_SUM_QTY_BUS_ADDR_WIDTH,
    INDEX_WIDTH => INDEX_WIDTH,
    TAG_WIDTH => TAG_WIDTH
  )
  PORT MAP(
    kernel_cmd_valid => l_sum_qty_cmd_accm_inst_kernel_cmd_valid,
    kernel_cmd_ready => l_sum_qty_cmd_accm_inst_kernel_cmd_ready,
    kernel_cmd_firstIdx => l_sum_qty_cmd_accm_inst_kernel_cmd_firstIdx,
    kernel_cmd_lastIdx => l_sum_qty_cmd_accm_inst_kernel_cmd_lastIdx,
    kernel_cmd_tag => l_sum_qty_cmd_accm_inst_kernel_cmd_tag,
    nucleus_cmd_valid => l_sum_qty_cmd_accm_inst_nucleus_cmd_valid,
    nucleus_cmd_ready => l_sum_qty_cmd_accm_inst_nucleus_cmd_ready,
    nucleus_cmd_firstIdx => l_sum_qty_cmd_accm_inst_nucleus_cmd_firstIdx,
    nucleus_cmd_lastIdx => l_sum_qty_cmd_accm_inst_nucleus_cmd_lastIdx,
    nucleus_cmd_ctrl => l_sum_qty_cmd_accm_inst_nucleus_cmd_ctrl,
    nucleus_cmd_tag => l_sum_qty_cmd_accm_inst_nucleus_cmd_tag,
    ctrl => l_sum_qty_cmd_accm_inst_ctrl
  );

  l_sum_base_price_cmd_accm_inst : ArrayCmdCtrlMerger
  GENERIC MAP(
    NUM_ADDR => 1,
    BUS_ADDR_WIDTH => L_SUM_BASE_PRICE_BUS_ADDR_WIDTH,
    INDEX_WIDTH => INDEX_WIDTH,
    TAG_WIDTH => TAG_WIDTH
  )
  PORT MAP(
    kernel_cmd_valid => l_sum_base_price_cmd_accm_inst_kernel_cmd_valid,
    kernel_cmd_ready => l_sum_base_price_cmd_accm_inst_kernel_cmd_ready,
    kernel_cmd_firstIdx => l_sum_base_price_cmd_accm_inst_kernel_cmd_firstIdx,
    kernel_cmd_lastIdx => l_sum_base_price_cmd_accm_inst_kernel_cmd_lastIdx,
    kernel_cmd_tag => l_sum_base_price_cmd_accm_inst_kernel_cmd_tag,
    nucleus_cmd_valid => l_sum_base_price_cmd_accm_inst_nucleus_cmd_valid,
    nucleus_cmd_ready => l_sum_base_price_cmd_accm_inst_nucleus_cmd_ready,
    nucleus_cmd_firstIdx => l_sum_base_price_cmd_accm_inst_nucleus_cmd_firstIdx,
    nucleus_cmd_lastIdx => l_sum_base_price_cmd_accm_inst_nucleus_cmd_lastIdx,
    nucleus_cmd_ctrl => l_sum_base_price_cmd_accm_inst_nucleus_cmd_ctrl,
    nucleus_cmd_tag => l_sum_base_price_cmd_accm_inst_nucleus_cmd_tag,
    ctrl => l_sum_base_price_cmd_accm_inst_ctrl
  );

  l_sum_disc_price_cmd_accm_inst : ArrayCmdCtrlMerger
  GENERIC MAP(
    NUM_ADDR => 1,
    BUS_ADDR_WIDTH => L_SUM_DISC_PRICE_BUS_ADDR_WIDTH,
    INDEX_WIDTH => INDEX_WIDTH,
    TAG_WIDTH => TAG_WIDTH
  )
  PORT MAP(
    kernel_cmd_valid => l_sum_disc_price_cmd_accm_inst_kernel_cmd_valid,
    kernel_cmd_ready => l_sum_disc_price_cmd_accm_inst_kernel_cmd_ready,
    kernel_cmd_firstIdx => l_sum_disc_price_cmd_accm_inst_kernel_cmd_firstIdx,
    kernel_cmd_lastIdx => l_sum_disc_price_cmd_accm_inst_kernel_cmd_lastIdx,
    kernel_cmd_tag => l_sum_disc_price_cmd_accm_inst_kernel_cmd_tag,
    nucleus_cmd_valid => l_sum_disc_price_cmd_accm_inst_nucleus_cmd_valid,
    nucleus_cmd_ready => l_sum_disc_price_cmd_accm_inst_nucleus_cmd_ready,
    nucleus_cmd_firstIdx => l_sum_disc_price_cmd_accm_inst_nucleus_cmd_firstIdx,
    nucleus_cmd_lastIdx => l_sum_disc_price_cmd_accm_inst_nucleus_cmd_lastIdx,
    nucleus_cmd_ctrl => l_sum_disc_price_cmd_accm_inst_nucleus_cmd_ctrl,
    nucleus_cmd_tag => l_sum_disc_price_cmd_accm_inst_nucleus_cmd_tag,
    ctrl => l_sum_disc_price_cmd_accm_inst_ctrl
  );

  l_sum_charge_cmd_accm_inst : ArrayCmdCtrlMerger
  GENERIC MAP(
    NUM_ADDR => 1,
    BUS_ADDR_WIDTH => L_SUM_CHARGE_BUS_ADDR_WIDTH,
    INDEX_WIDTH => INDEX_WIDTH,
    TAG_WIDTH => TAG_WIDTH
  )
  PORT MAP(
    kernel_cmd_valid => l_sum_charge_cmd_accm_inst_kernel_cmd_valid,
    kernel_cmd_ready => l_sum_charge_cmd_accm_inst_kernel_cmd_ready,
    kernel_cmd_firstIdx => l_sum_charge_cmd_accm_inst_kernel_cmd_firstIdx,
    kernel_cmd_lastIdx => l_sum_charge_cmd_accm_inst_kernel_cmd_lastIdx,
    kernel_cmd_tag => l_sum_charge_cmd_accm_inst_kernel_cmd_tag,
    nucleus_cmd_valid => l_sum_charge_cmd_accm_inst_nucleus_cmd_valid,
    nucleus_cmd_ready => l_sum_charge_cmd_accm_inst_nucleus_cmd_ready,
    nucleus_cmd_firstIdx => l_sum_charge_cmd_accm_inst_nucleus_cmd_firstIdx,
    nucleus_cmd_lastIdx => l_sum_charge_cmd_accm_inst_nucleus_cmd_lastIdx,
    nucleus_cmd_ctrl => l_sum_charge_cmd_accm_inst_nucleus_cmd_ctrl,
    nucleus_cmd_tag => l_sum_charge_cmd_accm_inst_nucleus_cmd_tag,
    ctrl => l_sum_charge_cmd_accm_inst_ctrl
  );

  l_avg_qty_cmd_accm_inst : ArrayCmdCtrlMerger
  GENERIC MAP(
    NUM_ADDR => 1,
    BUS_ADDR_WIDTH => L_AVG_QTY_BUS_ADDR_WIDTH,
    INDEX_WIDTH => INDEX_WIDTH,
    TAG_WIDTH => TAG_WIDTH
  )
  PORT MAP(
    kernel_cmd_valid => l_avg_qty_cmd_accm_inst_kernel_cmd_valid,
    kernel_cmd_ready => l_avg_qty_cmd_accm_inst_kernel_cmd_ready,
    kernel_cmd_firstIdx => l_avg_qty_cmd_accm_inst_kernel_cmd_firstIdx,
    kernel_cmd_lastIdx => l_avg_qty_cmd_accm_inst_kernel_cmd_lastIdx,
    kernel_cmd_tag => l_avg_qty_cmd_accm_inst_kernel_cmd_tag,
    nucleus_cmd_valid => l_avg_qty_cmd_accm_inst_nucleus_cmd_valid,
    nucleus_cmd_ready => l_avg_qty_cmd_accm_inst_nucleus_cmd_ready,
    nucleus_cmd_firstIdx => l_avg_qty_cmd_accm_inst_nucleus_cmd_firstIdx,
    nucleus_cmd_lastIdx => l_avg_qty_cmd_accm_inst_nucleus_cmd_lastIdx,
    nucleus_cmd_ctrl => l_avg_qty_cmd_accm_inst_nucleus_cmd_ctrl,
    nucleus_cmd_tag => l_avg_qty_cmd_accm_inst_nucleus_cmd_tag,
    ctrl => l_avg_qty_cmd_accm_inst_ctrl
  );

  l_avg_price_cmd_accm_inst : ArrayCmdCtrlMerger
  GENERIC MAP(
    NUM_ADDR => 1,
    BUS_ADDR_WIDTH => L_AVG_PRICE_BUS_ADDR_WIDTH,
    INDEX_WIDTH => INDEX_WIDTH,
    TAG_WIDTH => TAG_WIDTH
  )
  PORT MAP(
    kernel_cmd_valid => l_avg_price_cmd_accm_inst_kernel_cmd_valid,
    kernel_cmd_ready => l_avg_price_cmd_accm_inst_kernel_cmd_ready,
    kernel_cmd_firstIdx => l_avg_price_cmd_accm_inst_kernel_cmd_firstIdx,
    kernel_cmd_lastIdx => l_avg_price_cmd_accm_inst_kernel_cmd_lastIdx,
    kernel_cmd_tag => l_avg_price_cmd_accm_inst_kernel_cmd_tag,
    nucleus_cmd_valid => l_avg_price_cmd_accm_inst_nucleus_cmd_valid,
    nucleus_cmd_ready => l_avg_price_cmd_accm_inst_nucleus_cmd_ready,
    nucleus_cmd_firstIdx => l_avg_price_cmd_accm_inst_nucleus_cmd_firstIdx,
    nucleus_cmd_lastIdx => l_avg_price_cmd_accm_inst_nucleus_cmd_lastIdx,
    nucleus_cmd_ctrl => l_avg_price_cmd_accm_inst_nucleus_cmd_ctrl,
    nucleus_cmd_tag => l_avg_price_cmd_accm_inst_nucleus_cmd_tag,
    ctrl => l_avg_price_cmd_accm_inst_ctrl
  );

  l_avg_disc_cmd_accm_inst : ArrayCmdCtrlMerger
  GENERIC MAP(
    NUM_ADDR => 1,
    BUS_ADDR_WIDTH => L_AVG_DISC_BUS_ADDR_WIDTH,
    INDEX_WIDTH => INDEX_WIDTH,
    TAG_WIDTH => TAG_WIDTH
  )
  PORT MAP(
    kernel_cmd_valid => l_avg_disc_cmd_accm_inst_kernel_cmd_valid,
    kernel_cmd_ready => l_avg_disc_cmd_accm_inst_kernel_cmd_ready,
    kernel_cmd_firstIdx => l_avg_disc_cmd_accm_inst_kernel_cmd_firstIdx,
    kernel_cmd_lastIdx => l_avg_disc_cmd_accm_inst_kernel_cmd_lastIdx,
    kernel_cmd_tag => l_avg_disc_cmd_accm_inst_kernel_cmd_tag,
    nucleus_cmd_valid => l_avg_disc_cmd_accm_inst_nucleus_cmd_valid,
    nucleus_cmd_ready => l_avg_disc_cmd_accm_inst_nucleus_cmd_ready,
    nucleus_cmd_firstIdx => l_avg_disc_cmd_accm_inst_nucleus_cmd_firstIdx,
    nucleus_cmd_lastIdx => l_avg_disc_cmd_accm_inst_nucleus_cmd_lastIdx,
    nucleus_cmd_ctrl => l_avg_disc_cmd_accm_inst_nucleus_cmd_ctrl,
    nucleus_cmd_tag => l_avg_disc_cmd_accm_inst_nucleus_cmd_tag,
    ctrl => l_avg_disc_cmd_accm_inst_ctrl
  );

  l_count_order_cmd_accm_inst : ArrayCmdCtrlMerger
  GENERIC MAP(
    NUM_ADDR => 1,
    BUS_ADDR_WIDTH => L_COUNT_ORDER_BUS_ADDR_WIDTH,
    INDEX_WIDTH => INDEX_WIDTH,
    TAG_WIDTH => TAG_WIDTH
  )
  PORT MAP(
    kernel_cmd_valid => l_count_order_cmd_accm_inst_kernel_cmd_valid,
    kernel_cmd_ready => l_count_order_cmd_accm_inst_kernel_cmd_ready,
    kernel_cmd_firstIdx => l_count_order_cmd_accm_inst_kernel_cmd_firstIdx,
    kernel_cmd_lastIdx => l_count_order_cmd_accm_inst_kernel_cmd_lastIdx,
    kernel_cmd_tag => l_count_order_cmd_accm_inst_kernel_cmd_tag,
    nucleus_cmd_valid => l_count_order_cmd_accm_inst_nucleus_cmd_valid,
    nucleus_cmd_ready => l_count_order_cmd_accm_inst_nucleus_cmd_ready,
    nucleus_cmd_firstIdx => l_count_order_cmd_accm_inst_nucleus_cmd_firstIdx,
    nucleus_cmd_lastIdx => l_count_order_cmd_accm_inst_nucleus_cmd_lastIdx,
    nucleus_cmd_ctrl => l_count_order_cmd_accm_inst_nucleus_cmd_ctrl,
    nucleus_cmd_tag => l_count_order_cmd_accm_inst_nucleus_cmd_tag,
    ctrl => l_count_order_cmd_accm_inst_ctrl
  );
  l_quantity_cmd_valid <= l_quantity_cmd_accm_inst_nucleus_cmd_valid;
  l_quantity_cmd_accm_inst_nucleus_cmd_ready <= l_quantity_cmd_ready;
  l_quantity_cmd_firstIdx <= l_quantity_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_quantity_cmd_lastIdx <= l_quantity_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_quantity_cmd_ctrl <= l_quantity_cmd_accm_inst_nucleus_cmd_ctrl;
  l_quantity_cmd_tag <= l_quantity_cmd_accm_inst_nucleus_cmd_tag;

  l_extendedprice_cmd_valid <= l_extendedprice_cmd_accm_inst_nucleus_cmd_valid;
  l_extendedprice_cmd_accm_inst_nucleus_cmd_ready <= l_extendedprice_cmd_ready;
  l_extendedprice_cmd_firstIdx <= l_extendedprice_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_extendedprice_cmd_lastIdx <= l_extendedprice_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_extendedprice_cmd_ctrl <= l_extendedprice_cmd_accm_inst_nucleus_cmd_ctrl;
  l_extendedprice_cmd_tag <= l_extendedprice_cmd_accm_inst_nucleus_cmd_tag;

  l_discount_cmd_valid <= l_discount_cmd_accm_inst_nucleus_cmd_valid;
  l_discount_cmd_accm_inst_nucleus_cmd_ready <= l_discount_cmd_ready;
  l_discount_cmd_firstIdx <= l_discount_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_discount_cmd_lastIdx <= l_discount_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_discount_cmd_ctrl <= l_discount_cmd_accm_inst_nucleus_cmd_ctrl;
  l_discount_cmd_tag <= l_discount_cmd_accm_inst_nucleus_cmd_tag;

  l_tax_cmd_valid <= l_tax_cmd_accm_inst_nucleus_cmd_valid;
  l_tax_cmd_accm_inst_nucleus_cmd_ready <= l_tax_cmd_ready;
  l_tax_cmd_firstIdx <= l_tax_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_tax_cmd_lastIdx <= l_tax_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_tax_cmd_ctrl <= l_tax_cmd_accm_inst_nucleus_cmd_ctrl;
  l_tax_cmd_tag <= l_tax_cmd_accm_inst_nucleus_cmd_tag;

  l_returnflag_cmd_valid <= l_returnflag_cmd_accm_inst_nucleus_cmd_valid;
  l_returnflag_cmd_accm_inst_nucleus_cmd_ready <= l_returnflag_cmd_ready;
  l_returnflag_cmd_firstIdx <= l_returnflag_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_returnflag_cmd_lastIdx <= l_returnflag_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_returnflag_cmd_ctrl <= l_returnflag_cmd_accm_inst_nucleus_cmd_ctrl;
  l_returnflag_cmd_tag <= l_returnflag_cmd_accm_inst_nucleus_cmd_tag;

  l_linestatus_cmd_valid <= l_linestatus_cmd_accm_inst_nucleus_cmd_valid;
  l_linestatus_cmd_accm_inst_nucleus_cmd_ready <= l_linestatus_cmd_ready;
  l_linestatus_cmd_firstIdx <= l_linestatus_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_linestatus_cmd_lastIdx <= l_linestatus_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_linestatus_cmd_ctrl <= l_linestatus_cmd_accm_inst_nucleus_cmd_ctrl;
  l_linestatus_cmd_tag <= l_linestatus_cmd_accm_inst_nucleus_cmd_tag;

  l_shipdate_cmd_valid <= l_shipdate_cmd_accm_inst_nucleus_cmd_valid;
  l_shipdate_cmd_accm_inst_nucleus_cmd_ready <= l_shipdate_cmd_ready;
  l_shipdate_cmd_firstIdx <= l_shipdate_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_shipdate_cmd_lastIdx <= l_shipdate_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_shipdate_cmd_ctrl <= l_shipdate_cmd_accm_inst_nucleus_cmd_ctrl;
  l_shipdate_cmd_tag <= l_shipdate_cmd_accm_inst_nucleus_cmd_tag;

  PriceSummary_inst_l_quantity_valid <= l_quantity_valid;
  l_quantity_ready <= PriceSummary_inst_l_quantity_ready;
  PriceSummary_inst_l_quantity_dvalid <= l_quantity_dvalid;
  PriceSummary_inst_l_quantity_last <= l_quantity_last;
  PriceSummary_inst_l_quantity <= l_quantity;

  PriceSummary_inst_l_extendedprice_valid <= l_extendedprice_valid;
  l_extendedprice_ready <= PriceSummary_inst_l_extendedprice_ready;
  PriceSummary_inst_l_extendedprice_dvalid <= l_extendedprice_dvalid;
  PriceSummary_inst_l_extendedprice_last <= l_extendedprice_last;
  PriceSummary_inst_l_extendedprice <= l_extendedprice;

  PriceSummary_inst_l_discount_valid <= l_discount_valid;
  l_discount_ready <= PriceSummary_inst_l_discount_ready;
  PriceSummary_inst_l_discount_dvalid <= l_discount_dvalid;
  PriceSummary_inst_l_discount_last <= l_discount_last;
  PriceSummary_inst_l_discount <= l_discount;

  PriceSummary_inst_l_tax_valid <= l_tax_valid;
  l_tax_ready <= PriceSummary_inst_l_tax_ready;
  PriceSummary_inst_l_tax_dvalid <= l_tax_dvalid;
  PriceSummary_inst_l_tax_last <= l_tax_last;
  PriceSummary_inst_l_tax <= l_tax;

  PriceSummary_inst_l_returnflag_valid <= l_returnflag_valid;
  l_returnflag_ready <= PriceSummary_inst_l_returnflag_ready;
  PriceSummary_inst_l_returnflag_dvalid <= l_returnflag_dvalid;
  PriceSummary_inst_l_returnflag_last <= l_returnflag_last;
  PriceSummary_inst_l_returnflag_length <= l_returnflag_length;
  PriceSummary_inst_l_returnflag_count <= l_returnflag_count;
  PriceSummary_inst_l_returnflag_chars_valid <= l_returnflag_chars_valid;
  l_returnflag_chars_ready <= PriceSummary_inst_l_returnflag_chars_ready;
  PriceSummary_inst_l_returnflag_chars_dvalid <= l_returnflag_chars_dvalid;
  PriceSummary_inst_l_returnflag_chars_last <= l_returnflag_chars_last;
  PriceSummary_inst_l_returnflag_chars <= l_returnflag_chars;
  PriceSummary_inst_l_returnflag_chars_count <= l_returnflag_chars_count;

  PriceSummary_inst_l_linestatus_valid <= l_linestatus_valid;
  l_linestatus_ready <= PriceSummary_inst_l_linestatus_ready;
  PriceSummary_inst_l_linestatus_dvalid <= l_linestatus_dvalid;
  PriceSummary_inst_l_linestatus_last <= l_linestatus_last;
  PriceSummary_inst_l_linestatus_length <= l_linestatus_length;
  PriceSummary_inst_l_linestatus_count <= l_linestatus_count;
  PriceSummary_inst_l_linestatus_chars_valid <= l_linestatus_chars_valid;
  l_linestatus_chars_ready <= PriceSummary_inst_l_linestatus_chars_ready;
  PriceSummary_inst_l_linestatus_chars_dvalid <= l_linestatus_chars_dvalid;
  PriceSummary_inst_l_linestatus_chars_last <= l_linestatus_chars_last;
  PriceSummary_inst_l_linestatus_chars <= l_linestatus_chars;
  PriceSummary_inst_l_linestatus_chars_count <= l_linestatus_chars_count;

  PriceSummary_inst_l_shipdate_valid <= l_shipdate_valid;
  l_shipdate_ready <= PriceSummary_inst_l_shipdate_ready;
  PriceSummary_inst_l_shipdate_dvalid <= l_shipdate_dvalid;
  PriceSummary_inst_l_shipdate_last <= l_shipdate_last;
  PriceSummary_inst_l_shipdate <= l_shipdate;

  PriceSummary_inst_l_quantity_unl_valid <= l_quantity_unl_valid;
  l_quantity_unl_ready <= PriceSummary_inst_l_quantity_unl_ready;
  PriceSummary_inst_l_quantity_unl_tag <= l_quantity_unl_tag;

  PriceSummary_inst_l_extendedprice_unl_valid <= l_extendedprice_unl_valid;
  l_extendedprice_unl_ready <= PriceSummary_inst_l_extendedprice_unl_ready;
  PriceSummary_inst_l_extendedprice_unl_tag <= l_extendedprice_unl_tag;

  PriceSummary_inst_l_discount_unl_valid <= l_discount_unl_valid;
  l_discount_unl_ready <= PriceSummary_inst_l_discount_unl_ready;
  PriceSummary_inst_l_discount_unl_tag <= l_discount_unl_tag;

  PriceSummary_inst_l_tax_unl_valid <= l_tax_unl_valid;
  l_tax_unl_ready <= PriceSummary_inst_l_tax_unl_ready;
  PriceSummary_inst_l_tax_unl_tag <= l_tax_unl_tag;

  PriceSummary_inst_l_returnflag_unl_valid <= l_returnflag_unl_valid;
  l_returnflag_unl_ready <= PriceSummary_inst_l_returnflag_unl_ready;
  PriceSummary_inst_l_returnflag_unl_tag <= l_returnflag_unl_tag;

  PriceSummary_inst_l_linestatus_unl_valid <= l_linestatus_unl_valid;
  l_linestatus_unl_ready <= PriceSummary_inst_l_linestatus_unl_ready;
  PriceSummary_inst_l_linestatus_unl_tag <= l_linestatus_unl_tag;

  PriceSummary_inst_l_shipdate_unl_valid <= l_shipdate_unl_valid;
  l_shipdate_unl_ready <= PriceSummary_inst_l_shipdate_unl_ready;
  PriceSummary_inst_l_shipdate_unl_tag <= l_shipdate_unl_tag;

  PriceSummary_inst_start <= mmio_inst_f_start_data;
  PriceSummary_inst_stop <= mmio_inst_f_stop_data;
  PriceSummary_inst_reset <= mmio_inst_f_reset_data;
  PriceSummary_inst_l_firstidx <= mmio_inst_f_l_firstidx_data;
  PriceSummary_inst_l_lastidx <= mmio_inst_f_l_lastidx_data;
  mmio_inst_f_idle_write_data <= PriceSummary_inst_idle;
  mmio_inst_f_busy_write_data <= PriceSummary_inst_busy;
  mmio_inst_f_done_write_data <= PriceSummary_inst_done;
  mmio_inst_f_result_write_data <= PriceSummary_inst_result;
  mmio_inst_f_rhigh_write_data <= PriceSummary_inst_rhigh;
  mmio_inst_f_rlow_write_data <= PriceSummary_inst_rlow;
  mmio_inst_f_status_1_write_data <= PriceSummary_inst_status_1;
  mmio_inst_f_status_2_write_data <= PriceSummary_inst_status_2;
  mmio_inst_f_r1_write_data <= PriceSummary_inst_r1;
  mmio_inst_f_r2_write_data <= PriceSummary_inst_r2;
  mmio_inst_f_r3_write_data <= PriceSummary_inst_r3;
  mmio_inst_f_r4_write_data <= PriceSummary_inst_r4;
  mmio_inst_f_r5_write_data <= PriceSummary_inst_r5;
  mmio_inst_f_r6_write_data <= PriceSummary_inst_r6;
  mmio_inst_f_r7_write_data <= PriceSummary_inst_r7;
  mmio_inst_f_r8_write_data <= PriceSummary_inst_r8;
  mmio_inst_mmio_awvalid <= mmio_awvalid;
  mmio_awready <= mmio_inst_mmio_awready;
  mmio_inst_mmio_awaddr <= mmio_awaddr;
  mmio_inst_mmio_wvalid <= mmio_wvalid;
  mmio_wready <= mmio_inst_mmio_wready;
  mmio_inst_mmio_wdata <= mmio_wdata;
  mmio_inst_mmio_wstrb <= mmio_wstrb;
  mmio_bvalid <= mmio_inst_mmio_bvalid;
  mmio_inst_mmio_bready <= mmio_bready;
  mmio_bresp <= mmio_inst_mmio_bresp;
  mmio_inst_mmio_arvalid <= mmio_arvalid;
  mmio_arready <= mmio_inst_mmio_arready;
  mmio_inst_mmio_araddr <= mmio_araddr;
  mmio_rvalid <= mmio_inst_mmio_rvalid;
  mmio_inst_mmio_rready <= mmio_rready;
  mmio_rdata <= mmio_inst_mmio_rdata;
  mmio_rresp <= mmio_inst_mmio_rresp;

  l_quantity_cmd_accm_inst_kernel_cmd_valid <= PriceSummary_inst_l_quantity_cmd_valid;
  PriceSummary_inst_l_quantity_cmd_ready <= l_quantity_cmd_accm_inst_kernel_cmd_ready;
  l_quantity_cmd_accm_inst_kernel_cmd_firstIdx <= PriceSummary_inst_l_quantity_cmd_firstIdx;
  l_quantity_cmd_accm_inst_kernel_cmd_lastIdx <= PriceSummary_inst_l_quantity_cmd_lastIdx;
  l_quantity_cmd_accm_inst_kernel_cmd_tag <= PriceSummary_inst_l_quantity_cmd_tag;

  l_extendedprice_cmd_accm_inst_kernel_cmd_valid <= PriceSummary_inst_l_extendedprice_cmd_valid;
  PriceSummary_inst_l_extendedprice_cmd_ready <= l_extendedprice_cmd_accm_inst_kernel_cmd_ready;
  l_extendedprice_cmd_accm_inst_kernel_cmd_firstIdx <= PriceSummary_inst_l_extendedprice_cmd_firstIdx;
  l_extendedprice_cmd_accm_inst_kernel_cmd_lastIdx <= PriceSummary_inst_l_extendedprice_cmd_lastIdx;
  l_extendedprice_cmd_accm_inst_kernel_cmd_tag <= PriceSummary_inst_l_extendedprice_cmd_tag;

  l_discount_cmd_accm_inst_kernel_cmd_valid <= PriceSummary_inst_l_discount_cmd_valid;
  PriceSummary_inst_l_discount_cmd_ready <= l_discount_cmd_accm_inst_kernel_cmd_ready;
  l_discount_cmd_accm_inst_kernel_cmd_firstIdx <= PriceSummary_inst_l_discount_cmd_firstIdx;
  l_discount_cmd_accm_inst_kernel_cmd_lastIdx <= PriceSummary_inst_l_discount_cmd_lastIdx;
  l_discount_cmd_accm_inst_kernel_cmd_tag <= PriceSummary_inst_l_discount_cmd_tag;

  l_tax_cmd_accm_inst_kernel_cmd_valid <= PriceSummary_inst_l_tax_cmd_valid;
  PriceSummary_inst_l_tax_cmd_ready <= l_tax_cmd_accm_inst_kernel_cmd_ready;
  l_tax_cmd_accm_inst_kernel_cmd_firstIdx <= PriceSummary_inst_l_tax_cmd_firstIdx;
  l_tax_cmd_accm_inst_kernel_cmd_lastIdx <= PriceSummary_inst_l_tax_cmd_lastIdx;
  l_tax_cmd_accm_inst_kernel_cmd_tag <= PriceSummary_inst_l_tax_cmd_tag;

  l_returnflag_cmd_accm_inst_kernel_cmd_valid <= PriceSummary_inst_l_returnflag_cmd_valid;
  PriceSummary_inst_l_returnflag_cmd_ready <= l_returnflag_cmd_accm_inst_kernel_cmd_ready;
  l_returnflag_cmd_accm_inst_kernel_cmd_firstIdx <= PriceSummary_inst_l_returnflag_cmd_firstIdx;
  l_returnflag_cmd_accm_inst_kernel_cmd_lastIdx <= PriceSummary_inst_l_returnflag_cmd_lastIdx;
  l_returnflag_cmd_accm_inst_kernel_cmd_tag <= PriceSummary_inst_l_returnflag_cmd_tag;

  l_linestatus_cmd_accm_inst_kernel_cmd_valid <= PriceSummary_inst_l_linestatus_cmd_valid;
  PriceSummary_inst_l_linestatus_cmd_ready <= l_linestatus_cmd_accm_inst_kernel_cmd_ready;
  l_linestatus_cmd_accm_inst_kernel_cmd_firstIdx <= PriceSummary_inst_l_linestatus_cmd_firstIdx;
  l_linestatus_cmd_accm_inst_kernel_cmd_lastIdx <= PriceSummary_inst_l_linestatus_cmd_lastIdx;
  l_linestatus_cmd_accm_inst_kernel_cmd_tag <= PriceSummary_inst_l_linestatus_cmd_tag;

  l_shipdate_cmd_accm_inst_kernel_cmd_valid <= PriceSummary_inst_l_shipdate_cmd_valid;
  PriceSummary_inst_l_shipdate_cmd_ready <= l_shipdate_cmd_accm_inst_kernel_cmd_ready;
  l_shipdate_cmd_accm_inst_kernel_cmd_firstIdx <= PriceSummary_inst_l_shipdate_cmd_firstIdx;
  l_shipdate_cmd_accm_inst_kernel_cmd_lastIdx <= PriceSummary_inst_l_shipdate_cmd_lastIdx;
  l_shipdate_cmd_accm_inst_kernel_cmd_tag <= PriceSummary_inst_l_shipdate_cmd_tag;

  l_quantity_cmd_accm_inst_ctrl(63 DOWNTO 0) <= mmio_inst_f_l_quantity_values_data;
  l_extendedprice_cmd_accm_inst_ctrl(63 DOWNTO 0) <= mmio_inst_f_l_extendedprice_values_data;
  l_discount_cmd_accm_inst_ctrl(63 DOWNTO 0) <= mmio_inst_f_l_discount_values_data;
  l_tax_cmd_accm_inst_ctrl(63 DOWNTO 0) <= mmio_inst_f_l_tax_values_data;
  l_returnflag_cmd_accm_inst_ctrl(63 DOWNTO 0) <= mmio_inst_f_l_returnflag_offsets_data;
  l_returnflag_cmd_accm_inst_ctrl(127 DOWNTO 64) <= mmio_inst_f_l_returnflag_values_data;

  l_linestatus_cmd_accm_inst_ctrl(63 DOWNTO 0) <= mmio_inst_f_l_linestatus_offsets_data;
  l_linestatus_cmd_accm_inst_ctrl(127 DOWNTO 64) <= mmio_inst_f_l_linestatus_values_data;

  l_shipdate_cmd_accm_inst_ctrl(63 DOWNTO 0) <= mmio_inst_f_l_shipdate_values_data;

  l_returnflag_o_valid <= PriceSummaryWriter_inst_l_returnflag_o_valid;
  PriceSummaryWriter_inst_l_returnflag_o_ready <= l_returnflag_o_ready;
  l_returnflag_o_dvalid <= PriceSummaryWriter_inst_l_returnflag_o_dvalid;
  l_returnflag_o_last <= PriceSummaryWriter_inst_l_returnflag_o_last;
  l_returnflag_o_length <= PriceSummaryWriter_inst_l_returnflag_o_length;
  l_returnflag_o_count <= PriceSummaryWriter_inst_l_returnflag_o_count;
  l_returnflag_o_chars_valid <= PriceSummaryWriter_inst_l_returnflag_o_chars_valid;
  PriceSummaryWriter_inst_l_returnflag_o_chars_ready <= l_returnflag_o_chars_ready;
  l_returnflag_o_chars_dvalid <= PriceSummaryWriter_inst_l_returnflag_o_chars_dvalid;
  l_returnflag_o_chars_last <= PriceSummaryWriter_inst_l_returnflag_o_chars_last;
  l_returnflag_o_chars <= PriceSummaryWriter_inst_l_returnflag_o_chars;
  l_returnflag_o_chars_count <= PriceSummaryWriter_inst_l_returnflag_o_chars_count;

  l_linestatus_o_valid <= PriceSummaryWriter_inst_l_linestatus_o_valid;
  PriceSummaryWriter_inst_l_linestatus_o_ready <= l_linestatus_o_ready;
  l_linestatus_o_dvalid <= PriceSummaryWriter_inst_l_linestatus_o_dvalid;
  l_linestatus_o_last <= PriceSummaryWriter_inst_l_linestatus_o_last;
  l_linestatus_o_length <= PriceSummaryWriter_inst_l_linestatus_o_length;
  l_linestatus_o_count <= PriceSummaryWriter_inst_l_linestatus_o_count;
  l_linestatus_o_chars_valid <= PriceSummaryWriter_inst_l_linestatus_o_chars_valid;
  PriceSummaryWriter_inst_l_linestatus_o_chars_ready <= l_linestatus_o_chars_ready;
  l_linestatus_o_chars_dvalid <= PriceSummaryWriter_inst_l_linestatus_o_chars_dvalid;
  l_linestatus_o_chars_last <= PriceSummaryWriter_inst_l_linestatus_o_chars_last;
  l_linestatus_o_chars <= PriceSummaryWriter_inst_l_linestatus_o_chars;
  l_linestatus_o_chars_count <= PriceSummaryWriter_inst_l_linestatus_o_chars_count;

  l_sum_qty_valid <= PriceSummaryWriter_inst_l_sum_qty_valid;
  PriceSummaryWriter_inst_l_sum_qty_ready <= l_sum_qty_ready;
  l_sum_qty_dvalid <= PriceSummaryWriter_inst_l_sum_qty_dvalid;
  l_sum_qty_last <= PriceSummaryWriter_inst_l_sum_qty_last;
  l_sum_qty <= PriceSummaryWriter_inst_l_sum_qty;

  l_sum_base_price_valid <= PriceSummaryWriter_inst_l_sum_base_price_valid;
  PriceSummaryWriter_inst_l_sum_base_price_ready <= l_sum_base_price_ready;
  l_sum_base_price_dvalid <= PriceSummaryWriter_inst_l_sum_base_price_dvalid;
  l_sum_base_price_last <= PriceSummaryWriter_inst_l_sum_base_price_last;
  l_sum_base_price <= PriceSummaryWriter_inst_l_sum_base_price;

  l_sum_disc_price_valid <= PriceSummaryWriter_inst_l_sum_disc_price_valid;
  PriceSummaryWriter_inst_l_sum_disc_price_ready <= l_sum_disc_price_ready;
  l_sum_disc_price_dvalid <= PriceSummaryWriter_inst_l_sum_disc_price_dvalid;
  l_sum_disc_price_last <= PriceSummaryWriter_inst_l_sum_disc_price_last;
  l_sum_disc_price <= PriceSummaryWriter_inst_l_sum_disc_price;

  l_sum_charge_valid <= PriceSummaryWriter_inst_l_sum_charge_valid;
  PriceSummaryWriter_inst_l_sum_charge_ready <= l_sum_charge_ready;
  l_sum_charge_dvalid <= PriceSummaryWriter_inst_l_sum_charge_dvalid;
  l_sum_charge_last <= PriceSummaryWriter_inst_l_sum_charge_last;
  l_sum_charge <= PriceSummaryWriter_inst_l_sum_charge;

  l_avg_qty_valid <= PriceSummaryWriter_inst_l_avg_qty_valid;
  PriceSummaryWriter_inst_l_avg_qty_ready <= l_avg_qty_ready;
  l_avg_qty_dvalid <= PriceSummaryWriter_inst_l_avg_qty_dvalid;
  l_avg_qty_last <= PriceSummaryWriter_inst_l_avg_qty_last;
  l_avg_qty <= PriceSummaryWriter_inst_l_avg_qty;

  l_avg_price_valid <= PriceSummaryWriter_inst_l_avg_price_valid;
  PriceSummaryWriter_inst_l_avg_price_ready <= l_avg_price_ready;
  l_avg_price_dvalid <= PriceSummaryWriter_inst_l_avg_price_dvalid;
  l_avg_price_last <= PriceSummaryWriter_inst_l_avg_price_last;
  l_avg_price <= PriceSummaryWriter_inst_l_avg_price;

  l_avg_disc_valid <= PriceSummaryWriter_inst_l_avg_disc_valid;
  PriceSummaryWriter_inst_l_avg_disc_ready <= l_avg_disc_ready;
  l_avg_disc_dvalid <= PriceSummaryWriter_inst_l_avg_disc_dvalid;
  l_avg_disc_last <= PriceSummaryWriter_inst_l_avg_disc_last;
  l_avg_disc <= PriceSummaryWriter_inst_l_avg_disc;

  l_count_order_valid <= PriceSummaryWriter_inst_l_count_order_valid;
  PriceSummaryWriter_inst_l_count_order_ready <= l_count_order_ready;
  l_count_order_dvalid <= PriceSummaryWriter_inst_l_count_order_dvalid;
  l_count_order_last <= PriceSummaryWriter_inst_l_count_order_last;
  l_count_order <= PriceSummaryWriter_inst_l_count_order;

  l_returnflag_o_cmd_valid <= l_returnflag_o_cmd_accm_inst_nucleus_cmd_valid;
  l_returnflag_o_cmd_accm_inst_nucleus_cmd_ready <= l_returnflag_o_cmd_ready;
  l_returnflag_o_cmd_firstIdx <= l_returnflag_o_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_returnflag_o_cmd_lastIdx <= l_returnflag_o_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_returnflag_o_cmd_ctrl <= l_returnflag_o_cmd_accm_inst_nucleus_cmd_ctrl;
  l_returnflag_o_cmd_tag <= l_returnflag_o_cmd_accm_inst_nucleus_cmd_tag;

  l_linestatus_o_cmd_valid <= l_linestatus_o_cmd_accm_inst_nucleus_cmd_valid;
  l_linestatus_o_cmd_accm_inst_nucleus_cmd_ready <= l_linestatus_o_cmd_ready;
  l_linestatus_o_cmd_firstIdx <= l_linestatus_o_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_linestatus_o_cmd_lastIdx <= l_linestatus_o_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_linestatus_o_cmd_ctrl <= l_linestatus_o_cmd_accm_inst_nucleus_cmd_ctrl;
  l_linestatus_o_cmd_tag <= l_linestatus_o_cmd_accm_inst_nucleus_cmd_tag;

  l_sum_qty_cmd_valid <= l_sum_qty_cmd_accm_inst_nucleus_cmd_valid;
  l_sum_qty_cmd_accm_inst_nucleus_cmd_ready <= l_sum_qty_cmd_ready;
  l_sum_qty_cmd_firstIdx <= l_sum_qty_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_sum_qty_cmd_lastIdx <= l_sum_qty_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_sum_qty_cmd_ctrl <= l_sum_qty_cmd_accm_inst_nucleus_cmd_ctrl;
  l_sum_qty_cmd_tag <= l_sum_qty_cmd_accm_inst_nucleus_cmd_tag;

  l_sum_base_price_cmd_valid <= l_sum_base_price_cmd_accm_inst_nucleus_cmd_valid;
  l_sum_base_price_cmd_accm_inst_nucleus_cmd_ready <= l_sum_base_price_cmd_ready;
  l_sum_base_price_cmd_firstIdx <= l_sum_base_price_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_sum_base_price_cmd_lastIdx <= l_sum_base_price_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_sum_base_price_cmd_ctrl <= l_sum_base_price_cmd_accm_inst_nucleus_cmd_ctrl;
  l_sum_base_price_cmd_tag <= l_sum_base_price_cmd_accm_inst_nucleus_cmd_tag;

  l_sum_disc_price_cmd_valid <= l_sum_disc_price_cmd_accm_inst_nucleus_cmd_valid;
  l_sum_disc_price_cmd_accm_inst_nucleus_cmd_ready <= l_sum_disc_price_cmd_ready;
  l_sum_disc_price_cmd_firstIdx <= l_sum_disc_price_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_sum_disc_price_cmd_lastIdx <= l_sum_disc_price_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_sum_disc_price_cmd_ctrl <= l_sum_disc_price_cmd_accm_inst_nucleus_cmd_ctrl;
  l_sum_disc_price_cmd_tag <= l_sum_disc_price_cmd_accm_inst_nucleus_cmd_tag;

  l_sum_charge_cmd_valid <= l_sum_charge_cmd_accm_inst_nucleus_cmd_valid;
  l_sum_charge_cmd_accm_inst_nucleus_cmd_ready <= l_sum_charge_cmd_ready;
  l_sum_charge_cmd_firstIdx <= l_sum_charge_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_sum_charge_cmd_lastIdx <= l_sum_charge_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_sum_charge_cmd_ctrl <= l_sum_charge_cmd_accm_inst_nucleus_cmd_ctrl;
  l_sum_charge_cmd_tag <= l_sum_charge_cmd_accm_inst_nucleus_cmd_tag;

  l_avg_qty_cmd_valid <= l_avg_qty_cmd_accm_inst_nucleus_cmd_valid;
  l_avg_qty_cmd_accm_inst_nucleus_cmd_ready <= l_avg_qty_cmd_ready;
  l_avg_qty_cmd_firstIdx <= l_avg_qty_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_avg_qty_cmd_lastIdx <= l_avg_qty_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_avg_qty_cmd_ctrl <= l_avg_qty_cmd_accm_inst_nucleus_cmd_ctrl;
  l_avg_qty_cmd_tag <= l_avg_qty_cmd_accm_inst_nucleus_cmd_tag;

  l_avg_price_cmd_valid <= l_avg_price_cmd_accm_inst_nucleus_cmd_valid;
  l_avg_price_cmd_accm_inst_nucleus_cmd_ready <= l_avg_price_cmd_ready;
  l_avg_price_cmd_firstIdx <= l_avg_price_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_avg_price_cmd_lastIdx <= l_avg_price_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_avg_price_cmd_ctrl <= l_avg_price_cmd_accm_inst_nucleus_cmd_ctrl;
  l_avg_price_cmd_tag <= l_avg_price_cmd_accm_inst_nucleus_cmd_tag;

  l_avg_disc_cmd_valid <= l_avg_disc_cmd_accm_inst_nucleus_cmd_valid;
  l_avg_disc_cmd_accm_inst_nucleus_cmd_ready <= l_avg_disc_cmd_ready;
  l_avg_disc_cmd_firstIdx <= l_avg_disc_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_avg_disc_cmd_lastIdx <= l_avg_disc_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_avg_disc_cmd_ctrl <= l_avg_disc_cmd_accm_inst_nucleus_cmd_ctrl;
  l_avg_disc_cmd_tag <= l_avg_disc_cmd_accm_inst_nucleus_cmd_tag;

  l_count_order_cmd_valid <= l_count_order_cmd_accm_inst_nucleus_cmd_valid;
  l_count_order_cmd_accm_inst_nucleus_cmd_ready <= l_count_order_cmd_ready;
  l_count_order_cmd_firstIdx <= l_count_order_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_count_order_cmd_lastIdx <= l_count_order_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_count_order_cmd_ctrl <= l_count_order_cmd_accm_inst_nucleus_cmd_ctrl;
  l_count_order_cmd_tag <= l_count_order_cmd_accm_inst_nucleus_cmd_tag;

  PriceSummaryWriter_inst_l_returnflag_o_unl_valid <= l_returnflag_o_unl_valid;
  l_returnflag_o_unl_ready <= PriceSummaryWriter_inst_l_returnflag_o_unl_ready;
  PriceSummaryWriter_inst_l_returnflag_o_unl_tag <= l_returnflag_o_unl_tag;

  PriceSummaryWriter_inst_l_linestatus_o_unl_valid <= l_linestatus_o_unl_valid;
  l_linestatus_o_unl_ready <= PriceSummaryWriter_inst_l_linestatus_o_unl_ready;
  PriceSummaryWriter_inst_l_linestatus_o_unl_tag <= l_linestatus_o_unl_tag;

  PriceSummaryWriter_inst_l_sum_qty_unl_valid <= l_sum_qty_unl_valid;
  l_sum_qty_unl_ready <= PriceSummaryWriter_inst_l_sum_qty_unl_ready;
  PriceSummaryWriter_inst_l_sum_qty_unl_tag <= l_sum_qty_unl_tag;

  PriceSummaryWriter_inst_l_sum_base_price_unl_valid <= l_sum_base_price_unl_valid;
  l_sum_base_price_unl_ready <= PriceSummaryWriter_inst_l_sum_base_price_unl_ready;
  PriceSummaryWriter_inst_l_sum_base_price_unl_tag <= l_sum_base_price_unl_tag;

  PriceSummaryWriter_inst_l_sum_disc_price_unl_valid <= l_sum_disc_price_unl_valid;
  l_sum_disc_price_unl_ready <= PriceSummaryWriter_inst_l_sum_disc_price_unl_ready;
  PriceSummaryWriter_inst_l_sum_disc_price_unl_tag <= l_sum_disc_price_unl_tag;

  PriceSummaryWriter_inst_l_sum_charge_unl_valid <= l_sum_charge_unl_valid;
  l_sum_charge_unl_ready <= PriceSummaryWriter_inst_l_sum_charge_unl_ready;
  PriceSummaryWriter_inst_l_sum_charge_unl_tag <= l_sum_charge_unl_tag;

  PriceSummaryWriter_inst_l_avg_qty_unl_valid <= l_avg_qty_unl_valid;
  l_avg_qty_unl_ready <= PriceSummaryWriter_inst_l_avg_qty_unl_ready;
  PriceSummaryWriter_inst_l_avg_qty_unl_tag <= l_avg_qty_unl_tag;

  PriceSummaryWriter_inst_l_avg_price_unl_valid <= l_avg_price_unl_valid;
  l_avg_price_unl_ready <= PriceSummaryWriter_inst_l_avg_price_unl_ready;
  PriceSummaryWriter_inst_l_avg_price_unl_tag <= l_avg_price_unl_tag;

  PriceSummaryWriter_inst_l_avg_disc_unl_valid <= l_avg_disc_unl_valid;
  l_avg_disc_unl_ready <= PriceSummaryWriter_inst_l_avg_disc_unl_ready;
  PriceSummaryWriter_inst_l_avg_disc_unl_tag <= l_avg_disc_unl_tag;

  PriceSummaryWriter_inst_l_count_order_unl_valid <= l_count_order_unl_valid;
  l_count_order_unl_ready <= PriceSummaryWriter_inst_l_count_order_unl_ready;
  PriceSummaryWriter_inst_l_count_order_unl_tag <= l_count_order_unl_tag;

  PriceSummaryWriter_inst_start <= mmio_inst_f_start_data;
  PriceSummaryWriter_inst_stop <= mmio_inst_f_stop_data;
  PriceSummaryWriter_inst_reset <= mmio_inst_f_reset_data;
  PriceSummaryWriter_inst_l_firstidx <= mmio_inst_f_l_firstidx_data;
  PriceSummaryWriter_inst_l_lastidx <= mmio_inst_f_l_lastidx_data;

  l_returnflag_o_cmd_accm_inst_kernel_cmd_valid <= PriceSummaryWriter_inst_l_returnflag_o_cmd_valid;
  PriceSummaryWriter_inst_l_returnflag_o_cmd_ready <= l_returnflag_o_cmd_accm_inst_kernel_cmd_ready;
  l_returnflag_o_cmd_accm_inst_kernel_cmd_firstIdx <= PriceSummaryWriter_inst_l_returnflag_o_cmd_firstIdx;
  l_returnflag_o_cmd_accm_inst_kernel_cmd_lastIdx <= PriceSummaryWriter_inst_l_returnflag_o_cmd_lastIdx;
  l_returnflag_o_cmd_accm_inst_kernel_cmd_tag <= PriceSummaryWriter_inst_l_returnflag_o_cmd_tag;

  l_linestatus_o_cmd_accm_inst_kernel_cmd_valid <= PriceSummaryWriter_inst_l_linestatus_o_cmd_valid;
  PriceSummaryWriter_inst_l_linestatus_o_cmd_ready <= l_linestatus_o_cmd_accm_inst_kernel_cmd_ready;
  l_linestatus_o_cmd_accm_inst_kernel_cmd_firstIdx <= PriceSummaryWriter_inst_l_linestatus_o_cmd_firstIdx;
  l_linestatus_o_cmd_accm_inst_kernel_cmd_lastIdx <= PriceSummaryWriter_inst_l_linestatus_o_cmd_lastIdx;
  l_linestatus_o_cmd_accm_inst_kernel_cmd_tag <= PriceSummaryWriter_inst_l_linestatus_o_cmd_tag;

  l_sum_qty_cmd_accm_inst_kernel_cmd_valid <= PriceSummaryWriter_inst_l_sum_qty_cmd_valid;
  PriceSummaryWriter_inst_l_sum_qty_cmd_ready <= l_sum_qty_cmd_accm_inst_kernel_cmd_ready;
  l_sum_qty_cmd_accm_inst_kernel_cmd_firstIdx <= PriceSummaryWriter_inst_l_sum_qty_cmd_firstIdx;
  l_sum_qty_cmd_accm_inst_kernel_cmd_lastIdx <= PriceSummaryWriter_inst_l_sum_qty_cmd_lastIdx;
  l_sum_qty_cmd_accm_inst_kernel_cmd_tag <= PriceSummaryWriter_inst_l_sum_qty_cmd_tag;

  l_sum_base_price_cmd_accm_inst_kernel_cmd_valid <= PriceSummaryWriter_inst_l_sum_base_price_cmd_valid;
  PriceSummaryWriter_inst_l_sum_base_price_cmd_ready <= l_sum_base_price_cmd_accm_inst_kernel_cmd_ready;
  l_sum_base_price_cmd_accm_inst_kernel_cmd_firstIdx <= PriceSummaryWriter_inst_l_sum_base_price_cmd_firstIdx;
  l_sum_base_price_cmd_accm_inst_kernel_cmd_lastIdx <= PriceSummaryWriter_inst_l_sum_base_price_cmd_lastIdx;
  l_sum_base_price_cmd_accm_inst_kernel_cmd_tag <= PriceSummaryWriter_inst_l_sum_base_price_cmd_tag;

  l_sum_disc_price_cmd_accm_inst_kernel_cmd_valid <= PriceSummaryWriter_inst_l_sum_disc_price_cmd_valid;
  PriceSummaryWriter_inst_l_sum_disc_price_cmd_ready <= l_sum_disc_price_cmd_accm_inst_kernel_cmd_ready;
  l_sum_disc_price_cmd_accm_inst_kernel_cmd_firstIdx <= PriceSummaryWriter_inst_l_sum_disc_price_cmd_firstIdx;
  l_sum_disc_price_cmd_accm_inst_kernel_cmd_lastIdx <= PriceSummaryWriter_inst_l_sum_disc_price_cmd_lastIdx;
  l_sum_disc_price_cmd_accm_inst_kernel_cmd_tag <= PriceSummaryWriter_inst_l_sum_disc_price_cmd_tag;

  l_sum_charge_cmd_accm_inst_kernel_cmd_valid <= PriceSummaryWriter_inst_l_sum_charge_cmd_valid;
  PriceSummaryWriter_inst_l_sum_charge_cmd_ready <= l_sum_charge_cmd_accm_inst_kernel_cmd_ready;
  l_sum_charge_cmd_accm_inst_kernel_cmd_firstIdx <= PriceSummaryWriter_inst_l_sum_charge_cmd_firstIdx;
  l_sum_charge_cmd_accm_inst_kernel_cmd_lastIdx <= PriceSummaryWriter_inst_l_sum_charge_cmd_lastIdx;
  l_sum_charge_cmd_accm_inst_kernel_cmd_tag <= PriceSummaryWriter_inst_l_sum_charge_cmd_tag;

  l_avg_qty_cmd_accm_inst_kernel_cmd_valid <= PriceSummaryWriter_inst_l_avg_qty_cmd_valid;
  PriceSummaryWriter_inst_l_avg_qty_cmd_ready <= l_avg_qty_cmd_accm_inst_kernel_cmd_ready;
  l_avg_qty_cmd_accm_inst_kernel_cmd_firstIdx <= PriceSummaryWriter_inst_l_avg_qty_cmd_firstIdx;
  l_avg_qty_cmd_accm_inst_kernel_cmd_lastIdx <= PriceSummaryWriter_inst_l_avg_qty_cmd_lastIdx;
  l_avg_qty_cmd_accm_inst_kernel_cmd_tag <= PriceSummaryWriter_inst_l_avg_qty_cmd_tag;

  l_avg_price_cmd_accm_inst_kernel_cmd_valid <= PriceSummaryWriter_inst_l_avg_price_cmd_valid;
  PriceSummaryWriter_inst_l_avg_price_cmd_ready <= l_avg_price_cmd_accm_inst_kernel_cmd_ready;
  l_avg_price_cmd_accm_inst_kernel_cmd_firstIdx <= PriceSummaryWriter_inst_l_avg_price_cmd_firstIdx;
  l_avg_price_cmd_accm_inst_kernel_cmd_lastIdx <= PriceSummaryWriter_inst_l_avg_price_cmd_lastIdx;
  l_avg_price_cmd_accm_inst_kernel_cmd_tag <= PriceSummaryWriter_inst_l_avg_price_cmd_tag;

  l_avg_disc_cmd_accm_inst_kernel_cmd_valid <= PriceSummaryWriter_inst_l_avg_disc_cmd_valid;
  PriceSummaryWriter_inst_l_avg_disc_cmd_ready <= l_avg_disc_cmd_accm_inst_kernel_cmd_ready;
  l_avg_disc_cmd_accm_inst_kernel_cmd_firstIdx <= PriceSummaryWriter_inst_l_avg_disc_cmd_firstIdx;
  l_avg_disc_cmd_accm_inst_kernel_cmd_lastIdx <= PriceSummaryWriter_inst_l_avg_disc_cmd_lastIdx;
  l_avg_disc_cmd_accm_inst_kernel_cmd_tag <= PriceSummaryWriter_inst_l_avg_disc_cmd_tag;

  l_count_order_cmd_accm_inst_kernel_cmd_valid <= PriceSummaryWriter_inst_l_count_order_cmd_valid;
  PriceSummaryWriter_inst_l_count_order_cmd_ready <= l_count_order_cmd_accm_inst_kernel_cmd_ready;
  l_count_order_cmd_accm_inst_kernel_cmd_firstIdx <= PriceSummaryWriter_inst_l_count_order_cmd_firstIdx;
  l_count_order_cmd_accm_inst_kernel_cmd_lastIdx <= PriceSummaryWriter_inst_l_count_order_cmd_lastIdx;
  l_count_order_cmd_accm_inst_kernel_cmd_tag <= PriceSummaryWriter_inst_l_count_order_cmd_tag;

  l_returnflag_o_cmd_accm_inst_ctrl(63 DOWNTO 0) <= mmio_inst_f_l_returnflag_o_offsets_data;
  l_returnflag_o_cmd_accm_inst_ctrl(127 DOWNTO 64) <= mmio_inst_f_l_returnflag_o_values_data;

  l_linestatus_o_cmd_accm_inst_ctrl(63 DOWNTO 0) <= mmio_inst_f_l_linestatus_o_offsets_data;
  l_linestatus_o_cmd_accm_inst_ctrl(127 DOWNTO 64) <= mmio_inst_f_l_linestatus_o_values_data;

  l_sum_qty_cmd_accm_inst_ctrl(63 DOWNTO 0) <= mmio_inst_f_l_sum_qty_values_data;
  l_sum_base_price_cmd_accm_inst_ctrl(63 DOWNTO 0) <= mmio_inst_f_l_sum_base_price_values_data;
  l_sum_disc_price_cmd_accm_inst_ctrl(63 DOWNTO 0) <= mmio_inst_f_l_sum_disc_price_values_data;
  l_sum_charge_cmd_accm_inst_ctrl(63 DOWNTO 0) <= mmio_inst_f_l_sum_charge_values_data;
  l_avg_qty_cmd_accm_inst_ctrl(63 DOWNTO 0) <= mmio_inst_f_l_avg_qty_values_data;
  l_avg_price_cmd_accm_inst_ctrl(63 DOWNTO 0) <= mmio_inst_f_l_avg_price_values_data;
  l_avg_disc_cmd_accm_inst_ctrl(63 DOWNTO 0) <= mmio_inst_f_l_avg_disc_values_data;
  l_count_order_cmd_accm_inst_ctrl(63 DOWNTO 0) <= mmio_inst_f_l_count_order_values_data;
END ARCHITECTURE;