-- Copyright 2018-2019 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
-- This file was generated by Fletchgen. Modify this file at your own risk.

LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.numeric_std.ALL;

LIBRARY work;
USE work.Interconnect_pkg.ALL;

ENTITY PriceSummary_Mantle IS
  GENERIC (
    INDEX_WIDTH : INTEGER := 32;
    TAG_WIDTH : INTEGER := 1;
    BUS_ADDR_WIDTH : INTEGER := 64;
    BUS_DATA_WIDTH : INTEGER := 512;
    BUS_LEN_WIDTH : INTEGER := 8;
    BUS_BURST_STEP_LEN : INTEGER := 1;
    BUS_BURST_MAX_LEN : INTEGER := 16
  );
  PORT (
    bcd_clk : IN STD_LOGIC;
    bcd_reset : IN STD_LOGIC;
    kcd_clk : IN STD_LOGIC;
    kcd_reset : IN STD_LOGIC;
    mmio_awvalid : IN STD_LOGIC;
    mmio_awready : OUT STD_LOGIC;
    mmio_awaddr : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    mmio_wvalid : IN STD_LOGIC;
    mmio_wready : OUT STD_LOGIC;
    mmio_wdata : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    mmio_wstrb : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
    mmio_bvalid : OUT STD_LOGIC;
    mmio_bready : IN STD_LOGIC;
    mmio_bresp : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    mmio_arvalid : IN STD_LOGIC;
    mmio_arready : OUT STD_LOGIC;
    mmio_araddr : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
    mmio_rvalid : OUT STD_LOGIC;
    mmio_rready : IN STD_LOGIC;
    mmio_rdata : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
    mmio_rresp : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
    rd_mst_rreq_valid : OUT STD_LOGIC;
    rd_mst_rreq_ready : IN STD_LOGIC;
    rd_mst_rreq_addr : OUT STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
    rd_mst_rreq_len : OUT STD_LOGIC_VECTOR(BUS_LEN_WIDTH - 1 DOWNTO 0);
    rd_mst_rdat_valid : IN STD_LOGIC;
    rd_mst_rdat_ready : OUT STD_LOGIC;
    rd_mst_rdat_data : IN STD_LOGIC_VECTOR(BUS_DATA_WIDTH - 1 DOWNTO 0);
    rd_mst_rdat_last : IN STD_LOGIC;
    wr_mst_wreq_valid : OUT STD_LOGIC;
    wr_mst_wreq_ready : IN STD_LOGIC;
    wr_mst_wreq_addr : OUT STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
    wr_mst_wreq_len : OUT STD_LOGIC_VECTOR(BUS_LEN_WIDTH - 1 DOWNTO 0);
    wr_mst_wdat_valid : OUT STD_LOGIC;
    wr_mst_wdat_ready : IN STD_LOGIC;
    wr_mst_wdat_data : OUT STD_LOGIC_VECTOR(BUS_DATA_WIDTH - 1 DOWNTO 0);
    wr_mst_wdat_strobe : OUT STD_LOGIC_VECTOR(BUS_DATA_WIDTH/8 - 1 DOWNTO 0);
    wr_mst_wdat_last : OUT STD_LOGIC
  );
END ENTITY;

ARCHITECTURE Implementation OF PriceSummary_Mantle IS
  COMPONENT PriceSummary_Nucleus IS
    GENERIC (
      INDEX_WIDTH : INTEGER := 32;
      TAG_WIDTH : INTEGER := 1;
      L_QUANTITY_BUS_ADDR_WIDTH : INTEGER := 64;
      L_EXTENDEDPRICE_BUS_ADDR_WIDTH : INTEGER := 64;
      L_DISCOUNT_BUS_ADDR_WIDTH : INTEGER := 64;
      L_TAX_BUS_ADDR_WIDTH : INTEGER := 64;
      L_RETURNFLAG_BUS_ADDR_WIDTH : INTEGER := 64;
      L_LINESTATUS_BUS_ADDR_WIDTH : INTEGER := 64;
      L_SHIPDATE_BUS_ADDR_WIDTH : INTEGER := 64;
      L_RETURNFLAG_O_BUS_ADDR_WIDTH : INTEGER := 64;
      L_LINESTATUS_O_BUS_ADDR_WIDTH : INTEGER := 64;
      L_SUM_QTY_BUS_ADDR_WIDTH : INTEGER := 64;
      L_SUM_BASE_PRICE_BUS_ADDR_WIDTH : INTEGER := 64;
      L_SUM_DISC_PRICE_BUS_ADDR_WIDTH : INTEGER := 64;
      L_SUM_CHARGE_BUS_ADDR_WIDTH : INTEGER := 64;
      L_AVG_QTY_BUS_ADDR_WIDTH : INTEGER := 64;
      L_AVG_PRICE_BUS_ADDR_WIDTH : INTEGER := 64;
      L_AVG_DISC_BUS_ADDR_WIDTH : INTEGER := 64;
      L_COUNT_ORDER_BUS_ADDR_WIDTH : INTEGER := 64
    );
    PORT (
      kcd_clk : IN STD_LOGIC;
      kcd_reset : IN STD_LOGIC;
      mmio_awvalid : IN STD_LOGIC;
      mmio_awready : OUT STD_LOGIC;
      mmio_awaddr : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      mmio_wvalid : IN STD_LOGIC;
      mmio_wready : OUT STD_LOGIC;
      mmio_wdata : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      mmio_wstrb : IN STD_LOGIC_VECTOR(3 DOWNTO 0);
      mmio_bvalid : OUT STD_LOGIC;
      mmio_bready : IN STD_LOGIC;
      mmio_bresp : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      mmio_arvalid : IN STD_LOGIC;
      mmio_arready : OUT STD_LOGIC;
      mmio_araddr : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      mmio_rvalid : OUT STD_LOGIC;
      mmio_rready : IN STD_LOGIC;
      mmio_rdata : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
      mmio_rresp : OUT STD_LOGIC_VECTOR(1 DOWNTO 0);
      l_quantity_valid : IN STD_LOGIC;
      l_quantity_ready : OUT STD_LOGIC;
      l_quantity_dvalid : IN STD_LOGIC;
      l_quantity_last : IN STD_LOGIC;
      l_quantity : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_extendedprice_valid : IN STD_LOGIC;
      l_extendedprice_ready : OUT STD_LOGIC;
      l_extendedprice_dvalid : IN STD_LOGIC;
      l_extendedprice_last : IN STD_LOGIC;
      l_extendedprice : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_discount_valid : IN STD_LOGIC;
      l_discount_ready : OUT STD_LOGIC;
      l_discount_dvalid : IN STD_LOGIC;
      l_discount_last : IN STD_LOGIC;
      l_discount : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_tax_valid : IN STD_LOGIC;
      l_tax_ready : OUT STD_LOGIC;
      l_tax_dvalid : IN STD_LOGIC;
      l_tax_last : IN STD_LOGIC;
      l_tax : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_returnflag_valid : IN STD_LOGIC;
      l_returnflag_ready : OUT STD_LOGIC;
      l_returnflag_dvalid : IN STD_LOGIC;
      l_returnflag_last : IN STD_LOGIC;
      l_returnflag_length : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      l_returnflag_count : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      l_returnflag_chars_valid : IN STD_LOGIC;
      l_returnflag_chars_ready : OUT STD_LOGIC;
      l_returnflag_chars_dvalid : IN STD_LOGIC;
      l_returnflag_chars_last : IN STD_LOGIC;
      l_returnflag_chars : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      l_returnflag_chars_count : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      l_linestatus_valid : IN STD_LOGIC;
      l_linestatus_ready : OUT STD_LOGIC;
      l_linestatus_dvalid : IN STD_LOGIC;
      l_linestatus_last : IN STD_LOGIC;
      l_linestatus_length : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      l_linestatus_count : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      l_linestatus_chars_valid : IN STD_LOGIC;
      l_linestatus_chars_ready : OUT STD_LOGIC;
      l_linestatus_chars_dvalid : IN STD_LOGIC;
      l_linestatus_chars_last : IN STD_LOGIC;
      l_linestatus_chars : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      l_linestatus_chars_count : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      l_shipdate_valid : IN STD_LOGIC;
      l_shipdate_ready : OUT STD_LOGIC;
      l_shipdate_dvalid : IN STD_LOGIC;
      l_shipdate_last : IN STD_LOGIC;
      l_shipdate : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      l_quantity_unl_valid : IN STD_LOGIC;
      l_quantity_unl_ready : OUT STD_LOGIC;
      l_quantity_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_extendedprice_unl_valid : IN STD_LOGIC;
      l_extendedprice_unl_ready : OUT STD_LOGIC;
      l_extendedprice_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_discount_unl_valid : IN STD_LOGIC;
      l_discount_unl_ready : OUT STD_LOGIC;
      l_discount_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_tax_unl_valid : IN STD_LOGIC;
      l_tax_unl_ready : OUT STD_LOGIC;
      l_tax_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_returnflag_unl_valid : IN STD_LOGIC;
      l_returnflag_unl_ready : OUT STD_LOGIC;
      l_returnflag_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_linestatus_unl_valid : IN STD_LOGIC;
      l_linestatus_unl_ready : OUT STD_LOGIC;
      l_linestatus_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_shipdate_unl_valid : IN STD_LOGIC;
      l_shipdate_unl_ready : OUT STD_LOGIC;
      l_shipdate_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_quantity_cmd_valid : OUT STD_LOGIC;
      l_quantity_cmd_ready : IN STD_LOGIC;
      l_quantity_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_quantity_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_quantity_cmd_ctrl : OUT STD_LOGIC_VECTOR(L_QUANTITY_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_quantity_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_extendedprice_cmd_valid : OUT STD_LOGIC;
      l_extendedprice_cmd_ready : IN STD_LOGIC;
      l_extendedprice_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_extendedprice_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_extendedprice_cmd_ctrl : OUT STD_LOGIC_VECTOR(L_EXTENDEDPRICE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_extendedprice_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_discount_cmd_valid : OUT STD_LOGIC;
      l_discount_cmd_ready : IN STD_LOGIC;
      l_discount_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_discount_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_discount_cmd_ctrl : OUT STD_LOGIC_VECTOR(L_DISCOUNT_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_discount_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_tax_cmd_valid : OUT STD_LOGIC;
      l_tax_cmd_ready : IN STD_LOGIC;
      l_tax_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_tax_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_tax_cmd_ctrl : OUT STD_LOGIC_VECTOR(L_TAX_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_tax_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_returnflag_cmd_valid : OUT STD_LOGIC;
      l_returnflag_cmd_ready : IN STD_LOGIC;
      l_returnflag_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_returnflag_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_returnflag_cmd_ctrl : OUT STD_LOGIC_VECTOR(L_RETURNFLAG_BUS_ADDR_WIDTH * 2 - 1 DOWNTO 0);
      l_returnflag_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_linestatus_cmd_valid : OUT STD_LOGIC;
      l_linestatus_cmd_ready : IN STD_LOGIC;
      l_linestatus_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_linestatus_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_linestatus_cmd_ctrl : OUT STD_LOGIC_VECTOR(L_LINESTATUS_BUS_ADDR_WIDTH * 2 - 1 DOWNTO 0);
      l_linestatus_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_shipdate_cmd_valid : OUT STD_LOGIC;
      l_shipdate_cmd_ready : IN STD_LOGIC;
      l_shipdate_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_shipdate_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_shipdate_cmd_ctrl : OUT STD_LOGIC_VECTOR(L_SHIPDATE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_shipdate_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_returnflag_o_valid : OUT STD_LOGIC;
      l_returnflag_o_ready : IN STD_LOGIC;
      l_returnflag_o_dvalid : OUT STD_LOGIC;
      l_returnflag_o_last : OUT STD_LOGIC;
      l_returnflag_o_length : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
      l_returnflag_o_count : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      l_returnflag_o_chars_valid : OUT STD_LOGIC;
      l_returnflag_o_chars_ready : IN STD_LOGIC;
      l_returnflag_o_chars_dvalid : OUT STD_LOGIC;
      l_returnflag_o_chars_last : OUT STD_LOGIC;
      l_returnflag_o_chars : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
      l_returnflag_o_chars_count : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      l_linestatus_o_valid : OUT STD_LOGIC;
      l_linestatus_o_ready : IN STD_LOGIC;
      l_linestatus_o_dvalid : OUT STD_LOGIC;
      l_linestatus_o_last : OUT STD_LOGIC;
      l_linestatus_o_length : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
      l_linestatus_o_count : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      l_linestatus_o_chars_valid : OUT STD_LOGIC;
      l_linestatus_o_chars_ready : IN STD_LOGIC;
      l_linestatus_o_chars_dvalid : OUT STD_LOGIC;
      l_linestatus_o_chars_last : OUT STD_LOGIC;
      l_linestatus_o_chars : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
      l_linestatus_o_chars_count : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      l_sum_qty_valid : OUT STD_LOGIC;
      l_sum_qty_ready : IN STD_LOGIC;
      l_sum_qty_dvalid : OUT STD_LOGIC;
      l_sum_qty_last : OUT STD_LOGIC;
      l_sum_qty : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_sum_base_price_valid : OUT STD_LOGIC;
      l_sum_base_price_ready : IN STD_LOGIC;
      l_sum_base_price_dvalid : OUT STD_LOGIC;
      l_sum_base_price_last : OUT STD_LOGIC;
      l_sum_base_price : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_sum_disc_price_valid : OUT STD_LOGIC;
      l_sum_disc_price_ready : IN STD_LOGIC;
      l_sum_disc_price_dvalid : OUT STD_LOGIC;
      l_sum_disc_price_last : OUT STD_LOGIC;
      l_sum_disc_price : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_sum_charge_valid : OUT STD_LOGIC;
      l_sum_charge_ready : IN STD_LOGIC;
      l_sum_charge_dvalid : OUT STD_LOGIC;
      l_sum_charge_last : OUT STD_LOGIC;
      l_sum_charge : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_avg_qty_valid : OUT STD_LOGIC;
      l_avg_qty_ready : IN STD_LOGIC;
      l_avg_qty_dvalid : OUT STD_LOGIC;
      l_avg_qty_last : OUT STD_LOGIC;
      l_avg_qty : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_avg_price_valid : OUT STD_LOGIC;
      l_avg_price_ready : IN STD_LOGIC;
      l_avg_price_dvalid : OUT STD_LOGIC;
      l_avg_price_last : OUT STD_LOGIC;
      l_avg_price : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_avg_disc_valid : OUT STD_LOGIC;
      l_avg_disc_ready : IN STD_LOGIC;
      l_avg_disc_dvalid : OUT STD_LOGIC;
      l_avg_disc_last : OUT STD_LOGIC;
      l_avg_disc : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_count_order_valid : OUT STD_LOGIC;
      l_count_order_ready : IN STD_LOGIC;
      l_count_order_dvalid : OUT STD_LOGIC;
      l_count_order_last : OUT STD_LOGIC;
      l_count_order : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_returnflag_o_unl_valid : IN STD_LOGIC;
      l_returnflag_o_unl_ready : OUT STD_LOGIC;
      l_returnflag_o_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_linestatus_o_unl_valid : IN STD_LOGIC;
      l_linestatus_o_unl_ready : OUT STD_LOGIC;
      l_linestatus_o_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_sum_qty_unl_valid : IN STD_LOGIC;
      l_sum_qty_unl_ready : OUT STD_LOGIC;
      l_sum_qty_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_sum_base_price_unl_valid : IN STD_LOGIC;
      l_sum_base_price_unl_ready : OUT STD_LOGIC;
      l_sum_base_price_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_sum_disc_price_unl_valid : IN STD_LOGIC;
      l_sum_disc_price_unl_ready : OUT STD_LOGIC;
      l_sum_disc_price_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_sum_charge_unl_valid : IN STD_LOGIC;
      l_sum_charge_unl_ready : OUT STD_LOGIC;
      l_sum_charge_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_avg_qty_unl_valid : IN STD_LOGIC;
      l_avg_qty_unl_ready : OUT STD_LOGIC;
      l_avg_qty_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_avg_price_unl_valid : IN STD_LOGIC;
      l_avg_price_unl_ready : OUT STD_LOGIC;
      l_avg_price_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_avg_disc_unl_valid : IN STD_LOGIC;
      l_avg_disc_unl_ready : OUT STD_LOGIC;
      l_avg_disc_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_count_order_unl_valid : IN STD_LOGIC;
      l_count_order_unl_ready : OUT STD_LOGIC;
      l_count_order_unl_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_returnflag_o_cmd_valid : OUT STD_LOGIC;
      l_returnflag_o_cmd_ready : IN STD_LOGIC;
      l_returnflag_o_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_returnflag_o_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_returnflag_o_cmd_ctrl : OUT STD_LOGIC_VECTOR(L_RETURNFLAG_O_BUS_ADDR_WIDTH * 2 - 1 DOWNTO 0);
      l_returnflag_o_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_linestatus_o_cmd_valid : OUT STD_LOGIC;
      l_linestatus_o_cmd_ready : IN STD_LOGIC;
      l_linestatus_o_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_linestatus_o_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_linestatus_o_cmd_ctrl : OUT STD_LOGIC_VECTOR(L_LINESTATUS_O_BUS_ADDR_WIDTH * 2 - 1 DOWNTO 0);
      l_linestatus_o_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_sum_qty_cmd_valid : OUT STD_LOGIC;
      l_sum_qty_cmd_ready : IN STD_LOGIC;
      l_sum_qty_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_sum_qty_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_sum_qty_cmd_ctrl : OUT STD_LOGIC_VECTOR(L_SUM_QTY_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_sum_qty_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_sum_base_price_cmd_valid : OUT STD_LOGIC;
      l_sum_base_price_cmd_ready : IN STD_LOGIC;
      l_sum_base_price_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_sum_base_price_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_sum_base_price_cmd_ctrl : OUT STD_LOGIC_VECTOR(L_SUM_BASE_PRICE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_sum_base_price_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_sum_disc_price_cmd_valid : OUT STD_LOGIC;
      l_sum_disc_price_cmd_ready : IN STD_LOGIC;
      l_sum_disc_price_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_sum_disc_price_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_sum_disc_price_cmd_ctrl : OUT STD_LOGIC_VECTOR(L_SUM_DISC_PRICE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_sum_disc_price_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_sum_charge_cmd_valid : OUT STD_LOGIC;
      l_sum_charge_cmd_ready : IN STD_LOGIC;
      l_sum_charge_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_sum_charge_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_sum_charge_cmd_ctrl : OUT STD_LOGIC_VECTOR(L_SUM_CHARGE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_sum_charge_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_avg_qty_cmd_valid : OUT STD_LOGIC;
      l_avg_qty_cmd_ready : IN STD_LOGIC;
      l_avg_qty_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_avg_qty_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_avg_qty_cmd_ctrl : OUT STD_LOGIC_VECTOR(L_AVG_QTY_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_avg_qty_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_avg_price_cmd_valid : OUT STD_LOGIC;
      l_avg_price_cmd_ready : IN STD_LOGIC;
      l_avg_price_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_avg_price_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_avg_price_cmd_ctrl : OUT STD_LOGIC_VECTOR(L_AVG_PRICE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_avg_price_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_avg_disc_cmd_valid : OUT STD_LOGIC;
      l_avg_disc_cmd_ready : IN STD_LOGIC;
      l_avg_disc_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_avg_disc_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_avg_disc_cmd_ctrl : OUT STD_LOGIC_VECTOR(L_AVG_DISC_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_avg_disc_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_count_order_cmd_valid : OUT STD_LOGIC;
      l_count_order_cmd_ready : IN STD_LOGIC;
      l_count_order_cmd_firstIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_count_order_cmd_lastIdx : OUT STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_count_order_cmd_ctrl : OUT STD_LOGIC_VECTOR(L_COUNT_ORDER_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_count_order_cmd_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0)

    );
  END COMPONENT;

  COMPONENT PriceSummary_l IS
    GENERIC (
      INDEX_WIDTH : INTEGER := 32;
      TAG_WIDTH : INTEGER := 1;
      L_QUANTITY_BUS_ADDR_WIDTH : INTEGER := 64;
      L_QUANTITY_BUS_DATA_WIDTH : INTEGER := 512;
      L_QUANTITY_BUS_LEN_WIDTH : INTEGER := 8;
      L_QUANTITY_BUS_BURST_STEP_LEN : INTEGER := 1;
      L_QUANTITY_BUS_BURST_MAX_LEN : INTEGER := 16;
      L_EXTENDEDPRICE_BUS_ADDR_WIDTH : INTEGER := 64;
      L_EXTENDEDPRICE_BUS_DATA_WIDTH : INTEGER := 512;
      L_EXTENDEDPRICE_BUS_LEN_WIDTH : INTEGER := 8;
      L_EXTENDEDPRICE_BUS_BURST_STEP_LEN : INTEGER := 1;
      L_EXTENDEDPRICE_BUS_BURST_MAX_LEN : INTEGER := 16;
      L_DISCOUNT_BUS_ADDR_WIDTH : INTEGER := 64;
      L_DISCOUNT_BUS_DATA_WIDTH : INTEGER := 512;
      L_DISCOUNT_BUS_LEN_WIDTH : INTEGER := 8;
      L_DISCOUNT_BUS_BURST_STEP_LEN : INTEGER := 1;
      L_DISCOUNT_BUS_BURST_MAX_LEN : INTEGER := 16;
      L_TAX_BUS_ADDR_WIDTH : INTEGER := 64;
      L_TAX_BUS_DATA_WIDTH : INTEGER := 512;
      L_TAX_BUS_LEN_WIDTH : INTEGER := 8;
      L_TAX_BUS_BURST_STEP_LEN : INTEGER := 1;
      L_TAX_BUS_BURST_MAX_LEN : INTEGER := 16;
      L_RETURNFLAG_BUS_ADDR_WIDTH : INTEGER := 64;
      L_RETURNFLAG_BUS_DATA_WIDTH : INTEGER := 512;
      L_RETURNFLAG_BUS_LEN_WIDTH : INTEGER := 8;
      L_RETURNFLAG_BUS_BURST_STEP_LEN : INTEGER := 1;
      L_RETURNFLAG_BUS_BURST_MAX_LEN : INTEGER := 16;
      L_LINESTATUS_BUS_ADDR_WIDTH : INTEGER := 64;
      L_LINESTATUS_BUS_DATA_WIDTH : INTEGER := 512;
      L_LINESTATUS_BUS_LEN_WIDTH : INTEGER := 8;
      L_LINESTATUS_BUS_BURST_STEP_LEN : INTEGER := 1;
      L_LINESTATUS_BUS_BURST_MAX_LEN : INTEGER := 16;
      L_SHIPDATE_BUS_ADDR_WIDTH : INTEGER := 64;
      L_SHIPDATE_BUS_DATA_WIDTH : INTEGER := 512;
      L_SHIPDATE_BUS_LEN_WIDTH : INTEGER := 8;
      L_SHIPDATE_BUS_BURST_STEP_LEN : INTEGER := 1;
      L_SHIPDATE_BUS_BURST_MAX_LEN : INTEGER := 16;
      L_RETURNFLAG_O_BUS_ADDR_WIDTH : INTEGER := 64;
      L_RETURNFLAG_O_BUS_DATA_WIDTH : INTEGER := 512;
      L_RETURNFLAG_O_BUS_LEN_WIDTH : INTEGER := 8;
      L_RETURNFLAG_O_BUS_BURST_STEP_LEN : INTEGER := 1;
      L_RETURNFLAG_O_BUS_BURST_MAX_LEN : INTEGER := 16;
      L_LINESTATUS_O_BUS_ADDR_WIDTH : INTEGER := 64;
      L_LINESTATUS_O_BUS_DATA_WIDTH : INTEGER := 512;
      L_LINESTATUS_O_BUS_LEN_WIDTH : INTEGER := 8;
      L_LINESTATUS_O_BUS_BURST_STEP_LEN : INTEGER := 1;
      L_LINESTATUS_O_BUS_BURST_MAX_LEN : INTEGER := 16;
      L_SUM_QTY_BUS_ADDR_WIDTH : INTEGER := 64;
      L_SUM_QTY_BUS_DATA_WIDTH : INTEGER := 512;
      L_SUM_QTY_BUS_LEN_WIDTH : INTEGER := 8;
      L_SUM_QTY_BUS_BURST_STEP_LEN : INTEGER := 1;
      L_SUM_QTY_BUS_BURST_MAX_LEN : INTEGER := 16;
      L_SUM_BASE_PRICE_BUS_ADDR_WIDTH : INTEGER := 64;
      L_SUM_BASE_PRICE_BUS_DATA_WIDTH : INTEGER := 512;
      L_SUM_BASE_PRICE_BUS_LEN_WIDTH : INTEGER := 8;
      L_SUM_BASE_PRICE_BUS_BURST_STEP_LEN : INTEGER := 1;
      L_SUM_BASE_PRICE_BUS_BURST_MAX_LEN : INTEGER := 16;
      L_SUM_DISC_PRICE_BUS_ADDR_WIDTH : INTEGER := 64;
      L_SUM_DISC_PRICE_BUS_DATA_WIDTH : INTEGER := 512;
      L_SUM_DISC_PRICE_BUS_LEN_WIDTH : INTEGER := 8;
      L_SUM_DISC_PRICE_BUS_BURST_STEP_LEN : INTEGER := 1;
      L_SUM_DISC_PRICE_BUS_BURST_MAX_LEN : INTEGER := 16;
      L_SUM_CHARGE_BUS_ADDR_WIDTH : INTEGER := 64;
      L_SUM_CHARGE_BUS_DATA_WIDTH : INTEGER := 512;
      L_SUM_CHARGE_BUS_LEN_WIDTH : INTEGER := 8;
      L_SUM_CHARGE_BUS_BURST_STEP_LEN : INTEGER := 1;
      L_SUM_CHARGE_BUS_BURST_MAX_LEN : INTEGER := 16;
      L_AVG_QTY_BUS_ADDR_WIDTH : INTEGER := 64;
      L_AVG_QTY_BUS_DATA_WIDTH : INTEGER := 512;
      L_AVG_QTY_BUS_LEN_WIDTH : INTEGER := 8;
      L_AVG_QTY_BUS_BURST_STEP_LEN : INTEGER := 1;
      L_AVG_QTY_BUS_BURST_MAX_LEN : INTEGER := 16;
      L_AVG_PRICE_BUS_ADDR_WIDTH : INTEGER := 64;
      L_AVG_PRICE_BUS_DATA_WIDTH : INTEGER := 512;
      L_AVG_PRICE_BUS_LEN_WIDTH : INTEGER := 8;
      L_AVG_PRICE_BUS_BURST_STEP_LEN : INTEGER := 1;
      L_AVG_PRICE_BUS_BURST_MAX_LEN : INTEGER := 16;
      L_AVG_DISC_BUS_ADDR_WIDTH : INTEGER := 64;
      L_AVG_DISC_BUS_DATA_WIDTH : INTEGER := 512;
      L_AVG_DISC_BUS_LEN_WIDTH : INTEGER := 8;
      L_AVG_DISC_BUS_BURST_STEP_LEN : INTEGER := 1;
      L_AVG_DISC_BUS_BURST_MAX_LEN : INTEGER := 16;
      L_COUNT_ORDER_BUS_ADDR_WIDTH : INTEGER := 64;
      L_COUNT_ORDER_BUS_DATA_WIDTH : INTEGER := 512;
      L_COUNT_ORDER_BUS_LEN_WIDTH : INTEGER := 8;
      L_COUNT_ORDER_BUS_BURST_STEP_LEN : INTEGER := 1;
      L_COUNT_ORDER_BUS_BURST_MAX_LEN : INTEGER := 16
    );
    PORT (
      bcd_clk : IN STD_LOGIC;
      bcd_reset : IN STD_LOGIC;
      kcd_clk : IN STD_LOGIC;
      kcd_reset : IN STD_LOGIC;
      l_quantity_valid : OUT STD_LOGIC;
      l_quantity_ready : IN STD_LOGIC;
      l_quantity_dvalid : OUT STD_LOGIC;
      l_quantity_last : OUT STD_LOGIC;
      l_quantity : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_quantity_bus_rreq_valid : OUT STD_LOGIC;
      l_quantity_bus_rreq_ready : IN STD_LOGIC;
      l_quantity_bus_rreq_addr : OUT STD_LOGIC_VECTOR(L_QUANTITY_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_quantity_bus_rreq_len : OUT STD_LOGIC_VECTOR(L_QUANTITY_BUS_LEN_WIDTH - 1 DOWNTO 0);
      l_quantity_bus_rdat_valid : IN STD_LOGIC;
      l_quantity_bus_rdat_ready : OUT STD_LOGIC;
      l_quantity_bus_rdat_data : IN STD_LOGIC_VECTOR(L_QUANTITY_BUS_DATA_WIDTH - 1 DOWNTO 0);
      l_quantity_bus_rdat_last : IN STD_LOGIC;
      l_quantity_cmd_valid : IN STD_LOGIC;
      l_quantity_cmd_ready : OUT STD_LOGIC;
      l_quantity_cmd_firstIdx : IN STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_quantity_cmd_lastIdx : IN STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_quantity_cmd_ctrl : IN STD_LOGIC_VECTOR(L_QUANTITY_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_quantity_cmd_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_quantity_unl_valid : OUT STD_LOGIC;
      l_quantity_unl_ready : IN STD_LOGIC;
      l_quantity_unl_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_extendedprice_valid : OUT STD_LOGIC;
      l_extendedprice_ready : IN STD_LOGIC;
      l_extendedprice_dvalid : OUT STD_LOGIC;
      l_extendedprice_last : OUT STD_LOGIC;
      l_extendedprice : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_extendedprice_bus_rreq_valid : OUT STD_LOGIC;
      l_extendedprice_bus_rreq_ready : IN STD_LOGIC;
      l_extendedprice_bus_rreq_addr : OUT STD_LOGIC_VECTOR(L_EXTENDEDPRICE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_extendedprice_bus_rreq_len : OUT STD_LOGIC_VECTOR(L_EXTENDEDPRICE_BUS_LEN_WIDTH - 1 DOWNTO 0);
      l_extendedprice_bus_rdat_valid : IN STD_LOGIC;
      l_extendedprice_bus_rdat_ready : OUT STD_LOGIC;
      l_extendedprice_bus_rdat_data : IN STD_LOGIC_VECTOR(L_EXTENDEDPRICE_BUS_DATA_WIDTH - 1 DOWNTO 0);
      l_extendedprice_bus_rdat_last : IN STD_LOGIC;
      l_extendedprice_cmd_valid : IN STD_LOGIC;
      l_extendedprice_cmd_ready : OUT STD_LOGIC;
      l_extendedprice_cmd_firstIdx : IN STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_extendedprice_cmd_lastIdx : IN STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_extendedprice_cmd_ctrl : IN STD_LOGIC_VECTOR(L_EXTENDEDPRICE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_extendedprice_cmd_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_extendedprice_unl_valid : OUT STD_LOGIC;
      l_extendedprice_unl_ready : IN STD_LOGIC;
      l_extendedprice_unl_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_discount_valid : OUT STD_LOGIC;
      l_discount_ready : IN STD_LOGIC;
      l_discount_dvalid : OUT STD_LOGIC;
      l_discount_last : OUT STD_LOGIC;
      l_discount : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_discount_bus_rreq_valid : OUT STD_LOGIC;
      l_discount_bus_rreq_ready : IN STD_LOGIC;
      l_discount_bus_rreq_addr : OUT STD_LOGIC_VECTOR(L_DISCOUNT_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_discount_bus_rreq_len : OUT STD_LOGIC_VECTOR(L_DISCOUNT_BUS_LEN_WIDTH - 1 DOWNTO 0);
      l_discount_bus_rdat_valid : IN STD_LOGIC;
      l_discount_bus_rdat_ready : OUT STD_LOGIC;
      l_discount_bus_rdat_data : IN STD_LOGIC_VECTOR(L_DISCOUNT_BUS_DATA_WIDTH - 1 DOWNTO 0);
      l_discount_bus_rdat_last : IN STD_LOGIC;
      l_discount_cmd_valid : IN STD_LOGIC;
      l_discount_cmd_ready : OUT STD_LOGIC;
      l_discount_cmd_firstIdx : IN STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_discount_cmd_lastIdx : IN STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_discount_cmd_ctrl : IN STD_LOGIC_VECTOR(L_DISCOUNT_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_discount_cmd_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_discount_unl_valid : OUT STD_LOGIC;
      l_discount_unl_ready : IN STD_LOGIC;
      l_discount_unl_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_tax_valid : OUT STD_LOGIC;
      l_tax_ready : IN STD_LOGIC;
      l_tax_dvalid : OUT STD_LOGIC;
      l_tax_last : OUT STD_LOGIC;
      l_tax : OUT STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_tax_bus_rreq_valid : OUT STD_LOGIC;
      l_tax_bus_rreq_ready : IN STD_LOGIC;
      l_tax_bus_rreq_addr : OUT STD_LOGIC_VECTOR(L_TAX_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_tax_bus_rreq_len : OUT STD_LOGIC_VECTOR(L_TAX_BUS_LEN_WIDTH - 1 DOWNTO 0);
      l_tax_bus_rdat_valid : IN STD_LOGIC;
      l_tax_bus_rdat_ready : OUT STD_LOGIC;
      l_tax_bus_rdat_data : IN STD_LOGIC_VECTOR(L_TAX_BUS_DATA_WIDTH - 1 DOWNTO 0);
      l_tax_bus_rdat_last : IN STD_LOGIC;
      l_tax_cmd_valid : IN STD_LOGIC;
      l_tax_cmd_ready : OUT STD_LOGIC;
      l_tax_cmd_firstIdx : IN STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_tax_cmd_lastIdx : IN STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_tax_cmd_ctrl : IN STD_LOGIC_VECTOR(L_TAX_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_tax_cmd_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_tax_unl_valid : OUT STD_LOGIC;
      l_tax_unl_ready : IN STD_LOGIC;
      l_tax_unl_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_returnflag_valid : OUT STD_LOGIC;
      l_returnflag_ready : IN STD_LOGIC;
      l_returnflag_dvalid : OUT STD_LOGIC;
      l_returnflag_last : OUT STD_LOGIC;
      l_returnflag_length : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
      l_returnflag_count : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      l_returnflag_chars_valid : OUT STD_LOGIC;
      l_returnflag_chars_ready : IN STD_LOGIC;
      l_returnflag_chars_dvalid : OUT STD_LOGIC;
      l_returnflag_chars_last : OUT STD_LOGIC;
      l_returnflag_chars : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
      l_returnflag_chars_count : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      l_returnflag_bus_rreq_valid : OUT STD_LOGIC;
      l_returnflag_bus_rreq_ready : IN STD_LOGIC;
      l_returnflag_bus_rreq_addr : OUT STD_LOGIC_VECTOR(L_RETURNFLAG_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_returnflag_bus_rreq_len : OUT STD_LOGIC_VECTOR(L_RETURNFLAG_BUS_LEN_WIDTH - 1 DOWNTO 0);
      l_returnflag_bus_rdat_valid : IN STD_LOGIC;
      l_returnflag_bus_rdat_ready : OUT STD_LOGIC;
      l_returnflag_bus_rdat_data : IN STD_LOGIC_VECTOR(L_RETURNFLAG_BUS_DATA_WIDTH - 1 DOWNTO 0);
      l_returnflag_bus_rdat_last : IN STD_LOGIC;
      l_returnflag_cmd_valid : IN STD_LOGIC;
      l_returnflag_cmd_ready : OUT STD_LOGIC;
      l_returnflag_cmd_firstIdx : IN STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_returnflag_cmd_lastIdx : IN STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_returnflag_cmd_ctrl : IN STD_LOGIC_VECTOR(L_RETURNFLAG_BUS_ADDR_WIDTH * 2 - 1 DOWNTO 0);
      l_returnflag_cmd_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_returnflag_unl_valid : OUT STD_LOGIC;
      l_returnflag_unl_ready : IN STD_LOGIC;
      l_returnflag_unl_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_linestatus_valid : OUT STD_LOGIC;
      l_linestatus_ready : IN STD_LOGIC;
      l_linestatus_dvalid : OUT STD_LOGIC;
      l_linestatus_last : OUT STD_LOGIC;
      l_linestatus_length : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
      l_linestatus_count : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      l_linestatus_chars_valid : OUT STD_LOGIC;
      l_linestatus_chars_ready : IN STD_LOGIC;
      l_linestatus_chars_dvalid : OUT STD_LOGIC;
      l_linestatus_chars_last : OUT STD_LOGIC;
      l_linestatus_chars : OUT STD_LOGIC_VECTOR(7 DOWNTO 0);
      l_linestatus_chars_count : OUT STD_LOGIC_VECTOR(0 DOWNTO 0);
      l_linestatus_bus_rreq_valid : OUT STD_LOGIC;
      l_linestatus_bus_rreq_ready : IN STD_LOGIC;
      l_linestatus_bus_rreq_addr : OUT STD_LOGIC_VECTOR(L_LINESTATUS_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_linestatus_bus_rreq_len : OUT STD_LOGIC_VECTOR(L_LINESTATUS_BUS_LEN_WIDTH - 1 DOWNTO 0);
      l_linestatus_bus_rdat_valid : IN STD_LOGIC;
      l_linestatus_bus_rdat_ready : OUT STD_LOGIC;
      l_linestatus_bus_rdat_data : IN STD_LOGIC_VECTOR(L_LINESTATUS_BUS_DATA_WIDTH - 1 DOWNTO 0);
      l_linestatus_bus_rdat_last : IN STD_LOGIC;
      l_linestatus_cmd_valid : IN STD_LOGIC;
      l_linestatus_cmd_ready : OUT STD_LOGIC;
      l_linestatus_cmd_firstIdx : IN STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_linestatus_cmd_lastIdx : IN STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_linestatus_cmd_ctrl : IN STD_LOGIC_VECTOR(L_LINESTATUS_BUS_ADDR_WIDTH * 2 - 1 DOWNTO 0);
      l_linestatus_cmd_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_linestatus_unl_valid : OUT STD_LOGIC;
      l_linestatus_unl_ready : IN STD_LOGIC;
      l_linestatus_unl_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_shipdate_valid : OUT STD_LOGIC;
      l_shipdate_ready : IN STD_LOGIC;
      l_shipdate_dvalid : OUT STD_LOGIC;
      l_shipdate_last : OUT STD_LOGIC;
      l_shipdate : OUT STD_LOGIC_VECTOR(31 DOWNTO 0);
      l_shipdate_bus_rreq_valid : OUT STD_LOGIC;
      l_shipdate_bus_rreq_ready : IN STD_LOGIC;
      l_shipdate_bus_rreq_addr : OUT STD_LOGIC_VECTOR(L_SHIPDATE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_shipdate_bus_rreq_len : OUT STD_LOGIC_VECTOR(L_SHIPDATE_BUS_LEN_WIDTH - 1 DOWNTO 0);
      l_shipdate_bus_rdat_valid : IN STD_LOGIC;
      l_shipdate_bus_rdat_ready : OUT STD_LOGIC;
      l_shipdate_bus_rdat_data : IN STD_LOGIC_VECTOR(L_SHIPDATE_BUS_DATA_WIDTH - 1 DOWNTO 0);
      l_shipdate_bus_rdat_last : IN STD_LOGIC;
      l_shipdate_cmd_valid : IN STD_LOGIC;
      l_shipdate_cmd_ready : OUT STD_LOGIC;
      l_shipdate_cmd_firstIdx : IN STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_shipdate_cmd_lastIdx : IN STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_shipdate_cmd_ctrl : IN STD_LOGIC_VECTOR(L_SHIPDATE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_shipdate_cmd_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_shipdate_unl_valid : OUT STD_LOGIC;
      l_shipdate_unl_ready : IN STD_LOGIC;
      l_shipdate_unl_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_returnflag_o_valid : IN STD_LOGIC;
      l_returnflag_o_ready : OUT STD_LOGIC;
      l_returnflag_o_dvalid : IN STD_LOGIC;
      l_returnflag_o_last : IN STD_LOGIC;
      l_returnflag_o_length : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      l_returnflag_o_count : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      l_returnflag_o_chars_valid : IN STD_LOGIC;
      l_returnflag_o_chars_ready : OUT STD_LOGIC;
      l_returnflag_o_chars_dvalid : IN STD_LOGIC;
      l_returnflag_o_chars_last : IN STD_LOGIC;
      l_returnflag_o_chars : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      l_returnflag_o_chars_count : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      l_returnflag_o_bus_wreq_valid : OUT STD_LOGIC;
      l_returnflag_o_bus_wreq_ready : IN STD_LOGIC;
      l_returnflag_o_bus_wreq_addr : OUT STD_LOGIC_VECTOR(L_RETURNFLAG_O_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_returnflag_o_bus_wreq_len : OUT STD_LOGIC_VECTOR(L_RETURNFLAG_O_BUS_LEN_WIDTH - 1 DOWNTO 0);
      l_returnflag_o_bus_wdat_valid : OUT STD_LOGIC;
      l_returnflag_o_bus_wdat_ready : IN STD_LOGIC;
      l_returnflag_o_bus_wdat_data : OUT STD_LOGIC_VECTOR(L_RETURNFLAG_O_BUS_DATA_WIDTH - 1 DOWNTO 0);
      l_returnflag_o_bus_wdat_strobe : OUT STD_LOGIC_VECTOR(L_RETURNFLAG_O_BUS_DATA_WIDTH/8 - 1 DOWNTO 0);
      l_returnflag_o_bus_wdat_last : OUT STD_LOGIC;
      l_returnflag_o_cmd_valid : IN STD_LOGIC;
      l_returnflag_o_cmd_ready : OUT STD_LOGIC;
      l_returnflag_o_cmd_firstIdx : IN STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_returnflag_o_cmd_lastIdx : IN STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_returnflag_o_cmd_ctrl : IN STD_LOGIC_VECTOR(L_RETURNFLAG_O_BUS_ADDR_WIDTH * 2 - 1 DOWNTO 0);
      l_returnflag_o_cmd_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_returnflag_o_unl_valid : OUT STD_LOGIC;
      l_returnflag_o_unl_ready : IN STD_LOGIC;
      l_returnflag_o_unl_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_linestatus_o_valid : IN STD_LOGIC;
      l_linestatus_o_ready : OUT STD_LOGIC;
      l_linestatus_o_dvalid : IN STD_LOGIC;
      l_linestatus_o_last : IN STD_LOGIC;
      l_linestatus_o_length : IN STD_LOGIC_VECTOR(31 DOWNTO 0);
      l_linestatus_o_count : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      l_linestatus_o_chars_valid : IN STD_LOGIC;
      l_linestatus_o_chars_ready : OUT STD_LOGIC;
      l_linestatus_o_chars_dvalid : IN STD_LOGIC;
      l_linestatus_o_chars_last : IN STD_LOGIC;
      l_linestatus_o_chars : IN STD_LOGIC_VECTOR(7 DOWNTO 0);
      l_linestatus_o_chars_count : IN STD_LOGIC_VECTOR(0 DOWNTO 0);
      l_linestatus_o_bus_wreq_valid : OUT STD_LOGIC;
      l_linestatus_o_bus_wreq_ready : IN STD_LOGIC;
      l_linestatus_o_bus_wreq_addr : OUT STD_LOGIC_VECTOR(L_LINESTATUS_O_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_linestatus_o_bus_wreq_len : OUT STD_LOGIC_VECTOR(L_LINESTATUS_O_BUS_LEN_WIDTH - 1 DOWNTO 0);
      l_linestatus_o_bus_wdat_valid : OUT STD_LOGIC;
      l_linestatus_o_bus_wdat_ready : IN STD_LOGIC;
      l_linestatus_o_bus_wdat_data : OUT STD_LOGIC_VECTOR(L_LINESTATUS_O_BUS_DATA_WIDTH - 1 DOWNTO 0);
      l_linestatus_o_bus_wdat_strobe : OUT STD_LOGIC_VECTOR(L_LINESTATUS_O_BUS_DATA_WIDTH/8 - 1 DOWNTO 0);
      l_linestatus_o_bus_wdat_last : OUT STD_LOGIC;
      l_linestatus_o_cmd_valid : IN STD_LOGIC;
      l_linestatus_o_cmd_ready : OUT STD_LOGIC;
      l_linestatus_o_cmd_firstIdx : IN STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_linestatus_o_cmd_lastIdx : IN STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_linestatus_o_cmd_ctrl : IN STD_LOGIC_VECTOR(L_LINESTATUS_O_BUS_ADDR_WIDTH * 2 - 1 DOWNTO 0);
      l_linestatus_o_cmd_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_linestatus_o_unl_valid : OUT STD_LOGIC;
      l_linestatus_o_unl_ready : IN STD_LOGIC;
      l_linestatus_o_unl_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_sum_qty_valid : IN STD_LOGIC;
      l_sum_qty_ready : OUT STD_LOGIC;
      l_sum_qty_dvalid : IN STD_LOGIC;
      l_sum_qty_last : IN STD_LOGIC;
      l_sum_qty : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_sum_qty_bus_wreq_valid : OUT STD_LOGIC;
      l_sum_qty_bus_wreq_ready : IN STD_LOGIC;
      l_sum_qty_bus_wreq_addr : OUT STD_LOGIC_VECTOR(L_SUM_QTY_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_sum_qty_bus_wreq_len : OUT STD_LOGIC_VECTOR(L_SUM_QTY_BUS_LEN_WIDTH - 1 DOWNTO 0);
      l_sum_qty_bus_wdat_valid : OUT STD_LOGIC;
      l_sum_qty_bus_wdat_ready : IN STD_LOGIC;
      l_sum_qty_bus_wdat_data : OUT STD_LOGIC_VECTOR(L_SUM_QTY_BUS_DATA_WIDTH - 1 DOWNTO 0);
      l_sum_qty_bus_wdat_strobe : OUT STD_LOGIC_VECTOR(L_SUM_QTY_BUS_DATA_WIDTH/8 - 1 DOWNTO 0);
      l_sum_qty_bus_wdat_last : OUT STD_LOGIC;
      l_sum_qty_cmd_valid : IN STD_LOGIC;
      l_sum_qty_cmd_ready : OUT STD_LOGIC;
      l_sum_qty_cmd_firstIdx : IN STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_sum_qty_cmd_lastIdx : IN STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_sum_qty_cmd_ctrl : IN STD_LOGIC_VECTOR(L_SUM_QTY_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_sum_qty_cmd_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_sum_qty_unl_valid : OUT STD_LOGIC;
      l_sum_qty_unl_ready : IN STD_LOGIC;
      l_sum_qty_unl_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_sum_base_price_valid : IN STD_LOGIC;
      l_sum_base_price_ready : OUT STD_LOGIC;
      l_sum_base_price_dvalid : IN STD_LOGIC;
      l_sum_base_price_last : IN STD_LOGIC;
      l_sum_base_price : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_sum_base_price_bus_wreq_valid : OUT STD_LOGIC;
      l_sum_base_price_bus_wreq_ready : IN STD_LOGIC;
      l_sum_base_price_bus_wreq_addr : OUT STD_LOGIC_VECTOR(L_SUM_BASE_PRICE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_sum_base_price_bus_wreq_len : OUT STD_LOGIC_VECTOR(L_SUM_BASE_PRICE_BUS_LEN_WIDTH - 1 DOWNTO 0);
      l_sum_base_price_bus_wdat_valid : OUT STD_LOGIC;
      l_sum_base_price_bus_wdat_ready : IN STD_LOGIC;
      l_sum_base_price_bus_wdat_data : OUT STD_LOGIC_VECTOR(L_SUM_BASE_PRICE_BUS_DATA_WIDTH - 1 DOWNTO 0);
      l_sum_base_price_bus_wdat_strobe : OUT STD_LOGIC_VECTOR(L_SUM_BASE_PRICE_BUS_DATA_WIDTH/8 - 1 DOWNTO 0);
      l_sum_base_price_bus_wdat_last : OUT STD_LOGIC;
      l_sum_base_price_cmd_valid : IN STD_LOGIC;
      l_sum_base_price_cmd_ready : OUT STD_LOGIC;
      l_sum_base_price_cmd_firstIdx : IN STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_sum_base_price_cmd_lastIdx : IN STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_sum_base_price_cmd_ctrl : IN STD_LOGIC_VECTOR(L_SUM_BASE_PRICE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_sum_base_price_cmd_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_sum_base_price_unl_valid : OUT STD_LOGIC;
      l_sum_base_price_unl_ready : IN STD_LOGIC;
      l_sum_base_price_unl_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_sum_disc_price_valid : IN STD_LOGIC;
      l_sum_disc_price_ready : OUT STD_LOGIC;
      l_sum_disc_price_dvalid : IN STD_LOGIC;
      l_sum_disc_price_last : IN STD_LOGIC;
      l_sum_disc_price : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_sum_disc_price_bus_wreq_valid : OUT STD_LOGIC;
      l_sum_disc_price_bus_wreq_ready : IN STD_LOGIC;
      l_sum_disc_price_bus_wreq_addr : OUT STD_LOGIC_VECTOR(L_SUM_DISC_PRICE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_sum_disc_price_bus_wreq_len : OUT STD_LOGIC_VECTOR(L_SUM_DISC_PRICE_BUS_LEN_WIDTH - 1 DOWNTO 0);
      l_sum_disc_price_bus_wdat_valid : OUT STD_LOGIC;
      l_sum_disc_price_bus_wdat_ready : IN STD_LOGIC;
      l_sum_disc_price_bus_wdat_data : OUT STD_LOGIC_VECTOR(L_SUM_DISC_PRICE_BUS_DATA_WIDTH - 1 DOWNTO 0);
      l_sum_disc_price_bus_wdat_strobe : OUT STD_LOGIC_VECTOR(L_SUM_DISC_PRICE_BUS_DATA_WIDTH/8 - 1 DOWNTO 0);
      l_sum_disc_price_bus_wdat_last : OUT STD_LOGIC;
      l_sum_disc_price_cmd_valid : IN STD_LOGIC;
      l_sum_disc_price_cmd_ready : OUT STD_LOGIC;
      l_sum_disc_price_cmd_firstIdx : IN STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_sum_disc_price_cmd_lastIdx : IN STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_sum_disc_price_cmd_ctrl : IN STD_LOGIC_VECTOR(L_SUM_DISC_PRICE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_sum_disc_price_cmd_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_sum_disc_price_unl_valid : OUT STD_LOGIC;
      l_sum_disc_price_unl_ready : IN STD_LOGIC;
      l_sum_disc_price_unl_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_sum_charge_valid : IN STD_LOGIC;
      l_sum_charge_ready : OUT STD_LOGIC;
      l_sum_charge_dvalid : IN STD_LOGIC;
      l_sum_charge_last : IN STD_LOGIC;
      l_sum_charge : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_sum_charge_bus_wreq_valid : OUT STD_LOGIC;
      l_sum_charge_bus_wreq_ready : IN STD_LOGIC;
      l_sum_charge_bus_wreq_addr : OUT STD_LOGIC_VECTOR(L_SUM_CHARGE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_sum_charge_bus_wreq_len : OUT STD_LOGIC_VECTOR(L_SUM_CHARGE_BUS_LEN_WIDTH - 1 DOWNTO 0);
      l_sum_charge_bus_wdat_valid : OUT STD_LOGIC;
      l_sum_charge_bus_wdat_ready : IN STD_LOGIC;
      l_sum_charge_bus_wdat_data : OUT STD_LOGIC_VECTOR(L_SUM_CHARGE_BUS_DATA_WIDTH - 1 DOWNTO 0);
      l_sum_charge_bus_wdat_strobe : OUT STD_LOGIC_VECTOR(L_SUM_CHARGE_BUS_DATA_WIDTH/8 - 1 DOWNTO 0);
      l_sum_charge_bus_wdat_last : OUT STD_LOGIC;
      l_sum_charge_cmd_valid : IN STD_LOGIC;
      l_sum_charge_cmd_ready : OUT STD_LOGIC;
      l_sum_charge_cmd_firstIdx : IN STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_sum_charge_cmd_lastIdx : IN STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_sum_charge_cmd_ctrl : IN STD_LOGIC_VECTOR(L_SUM_CHARGE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_sum_charge_cmd_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_sum_charge_unl_valid : OUT STD_LOGIC;
      l_sum_charge_unl_ready : IN STD_LOGIC;
      l_sum_charge_unl_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_avg_qty_valid : IN STD_LOGIC;
      l_avg_qty_ready : OUT STD_LOGIC;
      l_avg_qty_dvalid : IN STD_LOGIC;
      l_avg_qty_last : IN STD_LOGIC;
      l_avg_qty : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_avg_qty_bus_wreq_valid : OUT STD_LOGIC;
      l_avg_qty_bus_wreq_ready : IN STD_LOGIC;
      l_avg_qty_bus_wreq_addr : OUT STD_LOGIC_VECTOR(L_AVG_QTY_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_avg_qty_bus_wreq_len : OUT STD_LOGIC_VECTOR(L_AVG_QTY_BUS_LEN_WIDTH - 1 DOWNTO 0);
      l_avg_qty_bus_wdat_valid : OUT STD_LOGIC;
      l_avg_qty_bus_wdat_ready : IN STD_LOGIC;
      l_avg_qty_bus_wdat_data : OUT STD_LOGIC_VECTOR(L_AVG_QTY_BUS_DATA_WIDTH - 1 DOWNTO 0);
      l_avg_qty_bus_wdat_strobe : OUT STD_LOGIC_VECTOR(L_AVG_QTY_BUS_DATA_WIDTH/8 - 1 DOWNTO 0);
      l_avg_qty_bus_wdat_last : OUT STD_LOGIC;
      l_avg_qty_cmd_valid : IN STD_LOGIC;
      l_avg_qty_cmd_ready : OUT STD_LOGIC;
      l_avg_qty_cmd_firstIdx : IN STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_avg_qty_cmd_lastIdx : IN STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_avg_qty_cmd_ctrl : IN STD_LOGIC_VECTOR(L_AVG_QTY_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_avg_qty_cmd_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_avg_qty_unl_valid : OUT STD_LOGIC;
      l_avg_qty_unl_ready : IN STD_LOGIC;
      l_avg_qty_unl_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_avg_price_valid : IN STD_LOGIC;
      l_avg_price_ready : OUT STD_LOGIC;
      l_avg_price_dvalid : IN STD_LOGIC;
      l_avg_price_last : IN STD_LOGIC;
      l_avg_price : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_avg_price_bus_wreq_valid : OUT STD_LOGIC;
      l_avg_price_bus_wreq_ready : IN STD_LOGIC;
      l_avg_price_bus_wreq_addr : OUT STD_LOGIC_VECTOR(L_AVG_PRICE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_avg_price_bus_wreq_len : OUT STD_LOGIC_VECTOR(L_AVG_PRICE_BUS_LEN_WIDTH - 1 DOWNTO 0);
      l_avg_price_bus_wdat_valid : OUT STD_LOGIC;
      l_avg_price_bus_wdat_ready : IN STD_LOGIC;
      l_avg_price_bus_wdat_data : OUT STD_LOGIC_VECTOR(L_AVG_PRICE_BUS_DATA_WIDTH - 1 DOWNTO 0);
      l_avg_price_bus_wdat_strobe : OUT STD_LOGIC_VECTOR(L_AVG_PRICE_BUS_DATA_WIDTH/8 - 1 DOWNTO 0);
      l_avg_price_bus_wdat_last : OUT STD_LOGIC;
      l_avg_price_cmd_valid : IN STD_LOGIC;
      l_avg_price_cmd_ready : OUT STD_LOGIC;
      l_avg_price_cmd_firstIdx : IN STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_avg_price_cmd_lastIdx : IN STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_avg_price_cmd_ctrl : IN STD_LOGIC_VECTOR(L_AVG_PRICE_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_avg_price_cmd_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_avg_price_unl_valid : OUT STD_LOGIC;
      l_avg_price_unl_ready : IN STD_LOGIC;
      l_avg_price_unl_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_avg_disc_valid : IN STD_LOGIC;
      l_avg_disc_ready : OUT STD_LOGIC;
      l_avg_disc_dvalid : IN STD_LOGIC;
      l_avg_disc_last : IN STD_LOGIC;
      l_avg_disc : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_avg_disc_bus_wreq_valid : OUT STD_LOGIC;
      l_avg_disc_bus_wreq_ready : IN STD_LOGIC;
      l_avg_disc_bus_wreq_addr : OUT STD_LOGIC_VECTOR(L_AVG_DISC_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_avg_disc_bus_wreq_len : OUT STD_LOGIC_VECTOR(L_AVG_DISC_BUS_LEN_WIDTH - 1 DOWNTO 0);
      l_avg_disc_bus_wdat_valid : OUT STD_LOGIC;
      l_avg_disc_bus_wdat_ready : IN STD_LOGIC;
      l_avg_disc_bus_wdat_data : OUT STD_LOGIC_VECTOR(L_AVG_DISC_BUS_DATA_WIDTH - 1 DOWNTO 0);
      l_avg_disc_bus_wdat_strobe : OUT STD_LOGIC_VECTOR(L_AVG_DISC_BUS_DATA_WIDTH/8 - 1 DOWNTO 0);
      l_avg_disc_bus_wdat_last : OUT STD_LOGIC;
      l_avg_disc_cmd_valid : IN STD_LOGIC;
      l_avg_disc_cmd_ready : OUT STD_LOGIC;
      l_avg_disc_cmd_firstIdx : IN STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_avg_disc_cmd_lastIdx : IN STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_avg_disc_cmd_ctrl : IN STD_LOGIC_VECTOR(L_AVG_DISC_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_avg_disc_cmd_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_avg_disc_unl_valid : OUT STD_LOGIC;
      l_avg_disc_unl_ready : IN STD_LOGIC;
      l_avg_disc_unl_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_count_order_valid : IN STD_LOGIC;
      l_count_order_ready : OUT STD_LOGIC;
      l_count_order_dvalid : IN STD_LOGIC;
      l_count_order_last : IN STD_LOGIC;
      l_count_order : IN STD_LOGIC_VECTOR(63 DOWNTO 0);
      l_count_order_bus_wreq_valid : OUT STD_LOGIC;
      l_count_order_bus_wreq_ready : IN STD_LOGIC;
      l_count_order_bus_wreq_addr : OUT STD_LOGIC_VECTOR(L_COUNT_ORDER_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_count_order_bus_wreq_len : OUT STD_LOGIC_VECTOR(L_COUNT_ORDER_BUS_LEN_WIDTH - 1 DOWNTO 0);
      l_count_order_bus_wdat_valid : OUT STD_LOGIC;
      l_count_order_bus_wdat_ready : IN STD_LOGIC;
      l_count_order_bus_wdat_data : OUT STD_LOGIC_VECTOR(L_COUNT_ORDER_BUS_DATA_WIDTH - 1 DOWNTO 0);
      l_count_order_bus_wdat_strobe : OUT STD_LOGIC_VECTOR(L_COUNT_ORDER_BUS_DATA_WIDTH/8 - 1 DOWNTO 0);
      l_count_order_bus_wdat_last : OUT STD_LOGIC;
      l_count_order_cmd_valid : IN STD_LOGIC;
      l_count_order_cmd_ready : OUT STD_LOGIC;
      l_count_order_cmd_firstIdx : IN STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_count_order_cmd_lastIdx : IN STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
      l_count_order_cmd_ctrl : IN STD_LOGIC_VECTOR(L_COUNT_ORDER_BUS_ADDR_WIDTH - 1 DOWNTO 0);
      l_count_order_cmd_tag : IN STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);
      l_count_order_unl_valid : OUT STD_LOGIC;
      l_count_order_unl_ready : IN STD_LOGIC;
      l_count_order_unl_tag : OUT STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0)
    );
  END COMPONENT;

  SIGNAL PriceSummaryWriter_Nucleus_inst_l_returnflag_o_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_returnflag_o_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_returnflag_o_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_returnflag_o_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_returnflag_o_length : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_returnflag_o_count : STD_LOGIC_VECTOR(0 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars : STD_LOGIC_VECTOR(7 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_count : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummaryWriter_Nucleus_inst_l_linestatus_o_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_linestatus_o_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_linestatus_o_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_linestatus_o_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_linestatus_o_length : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_linestatus_o_count : STD_LOGIC_VECTOR(0 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars : STD_LOGIC_VECTOR(7 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_count : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_qty_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_qty_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_qty_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_qty_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_qty : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_base_price_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_base_price_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_base_price_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_base_price_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_base_price : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_disc_price : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_charge_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_charge_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_charge_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_charge_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_charge : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_qty_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_qty_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_qty_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_qty_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_qty : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_price_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_price_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_price_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_price_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_price : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_disc_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_disc_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_disc_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_disc_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_disc : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummaryWriter_Nucleus_inst_l_count_order_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_count_order_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_count_order_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_count_order_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_count_order : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummaryWriter_Nucleus_inst_l_returnflag_o_unl_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_returnflag_o_unl_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_returnflag_o_unl_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_Nucleus_inst_l_linestatus_o_unl_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_linestatus_o_unl_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_linestatus_o_unl_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_qty_unl_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_qty_unl_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_qty_unl_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_base_price_unl_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_base_price_unl_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_base_price_unl_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_unl_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_unl_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_unl_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_charge_unl_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_charge_unl_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_charge_unl_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_qty_unl_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_qty_unl_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_qty_unl_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_price_unl_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_price_unl_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_price_unl_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_disc_unl_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_disc_unl_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_disc_unl_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_Nucleus_inst_l_count_order_unl_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_count_order_unl_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_count_order_unl_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_ctrl : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH * 2 - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_ctrl : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH * 2 - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_ctrl : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_ctrl : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_ctrl : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_ctrl : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_ctrl : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_ctrl : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_ctrl : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_ctrl : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_l_inst_l_returnflag_o_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_returnflag_o_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_returnflag_o_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_returnflag_o_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_returnflag_o_length : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_returnflag_o_count : STD_LOGIC_VECTOR(0 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_returnflag_o_chars_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_returnflag_o_chars_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_returnflag_o_chars_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_returnflag_o_chars_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_returnflag_o_chars : STD_LOGIC_VECTOR(7 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_returnflag_o_chars_count : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_addr : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_len : STD_LOGIC_VECTOR(BUS_LEN_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_data : STD_LOGIC_VECTOR(BUS_DATA_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_strobe : STD_LOGIC_VECTOR(BUS_DATA_WIDTH/8 - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_last : STD_LOGIC;

  SIGNAL PriceSummaryWriter_l_inst_l_returnflag_o_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_returnflag_o_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_returnflag_o_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_returnflag_o_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_returnflag_o_cmd_ctrl : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH * 2 - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_returnflag_o_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_l_inst_l_returnflag_o_unl_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_returnflag_o_unl_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_returnflag_o_unl_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_l_inst_l_linestatus_o_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_linestatus_o_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_linestatus_o_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_linestatus_o_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_linestatus_o_length : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_linestatus_o_count : STD_LOGIC_VECTOR(0 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_linestatus_o_chars_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_linestatus_o_chars_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_linestatus_o_chars_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_linestatus_o_chars_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_linestatus_o_chars : STD_LOGIC_VECTOR(7 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_linestatus_o_chars_count : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_addr : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_len : STD_LOGIC_VECTOR(BUS_LEN_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_data : STD_LOGIC_VECTOR(BUS_DATA_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_strobe : STD_LOGIC_VECTOR(BUS_DATA_WIDTH/8 - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_last : STD_LOGIC;

  SIGNAL PriceSummaryWriter_l_inst_l_linestatus_o_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_linestatus_o_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_linestatus_o_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_linestatus_o_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_linestatus_o_cmd_ctrl : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH * 2 - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_linestatus_o_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_l_inst_l_linestatus_o_unl_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_linestatus_o_unl_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_linestatus_o_unl_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_l_inst_l_sum_qty_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_qty_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_qty_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_qty_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_qty : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_addr : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_len : STD_LOGIC_VECTOR(BUS_LEN_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_data : STD_LOGIC_VECTOR(BUS_DATA_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_strobe : STD_LOGIC_VECTOR(BUS_DATA_WIDTH/8 - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_last : STD_LOGIC;

  SIGNAL PriceSummaryWriter_l_inst_l_sum_qty_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_qty_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_qty_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_sum_qty_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_sum_qty_cmd_ctrl : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_sum_qty_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_l_inst_l_sum_qty_unl_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_qty_unl_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_qty_unl_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_l_inst_l_sum_base_price_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_base_price_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_base_price_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_base_price_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_base_price : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_addr : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_len : STD_LOGIC_VECTOR(BUS_LEN_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_data : STD_LOGIC_VECTOR(BUS_DATA_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_strobe : STD_LOGIC_VECTOR(BUS_DATA_WIDTH/8 - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_last : STD_LOGIC;

  SIGNAL PriceSummaryWriter_l_inst_l_sum_base_price_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_base_price_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_base_price_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_sum_base_price_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_sum_base_price_cmd_ctrl : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_sum_base_price_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_l_inst_l_sum_base_price_unl_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_base_price_unl_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_base_price_unl_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_l_inst_l_sum_disc_price_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_disc_price_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_disc_price_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_disc_price_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_disc_price : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_addr : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_len : STD_LOGIC_VECTOR(BUS_LEN_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_data : STD_LOGIC_VECTOR(BUS_DATA_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_strobe : STD_LOGIC_VECTOR(BUS_DATA_WIDTH/8 - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_last : STD_LOGIC;

  SIGNAL PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_ctrl : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_l_inst_l_sum_disc_price_unl_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_disc_price_unl_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_disc_price_unl_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_l_inst_l_sum_charge_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_charge_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_charge_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_charge_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_charge : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_addr : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_len : STD_LOGIC_VECTOR(BUS_LEN_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_data : STD_LOGIC_VECTOR(BUS_DATA_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_strobe : STD_LOGIC_VECTOR(BUS_DATA_WIDTH/8 - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_last : STD_LOGIC;

  SIGNAL PriceSummaryWriter_l_inst_l_sum_charge_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_charge_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_charge_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_sum_charge_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_sum_charge_cmd_ctrl : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_sum_charge_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_l_inst_l_sum_charge_unl_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_charge_unl_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_sum_charge_unl_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_l_inst_l_avg_qty_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_qty_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_qty_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_qty_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_qty : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_addr : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_len : STD_LOGIC_VECTOR(BUS_LEN_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_data : STD_LOGIC_VECTOR(BUS_DATA_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_strobe : STD_LOGIC_VECTOR(BUS_DATA_WIDTH/8 - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_last : STD_LOGIC;

  SIGNAL PriceSummaryWriter_l_inst_l_avg_qty_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_qty_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_qty_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_avg_qty_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_avg_qty_cmd_ctrl : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_avg_qty_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_l_inst_l_avg_qty_unl_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_qty_unl_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_qty_unl_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_l_inst_l_avg_price_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_price_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_price_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_price_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_price : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_addr : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_len : STD_LOGIC_VECTOR(BUS_LEN_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_data : STD_LOGIC_VECTOR(BUS_DATA_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_strobe : STD_LOGIC_VECTOR(BUS_DATA_WIDTH/8 - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_last : STD_LOGIC;

  SIGNAL PriceSummaryWriter_l_inst_l_avg_price_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_price_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_price_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_avg_price_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_avg_price_cmd_ctrl : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_avg_price_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_l_inst_l_avg_price_unl_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_price_unl_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_price_unl_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_l_inst_l_avg_disc_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_disc_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_disc_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_disc_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_disc : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_addr : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_len : STD_LOGIC_VECTOR(BUS_LEN_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_data : STD_LOGIC_VECTOR(BUS_DATA_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_strobe : STD_LOGIC_VECTOR(BUS_DATA_WIDTH/8 - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_last : STD_LOGIC;

  SIGNAL PriceSummaryWriter_l_inst_l_avg_disc_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_disc_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_disc_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_avg_disc_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_avg_disc_cmd_ctrl : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_avg_disc_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_l_inst_l_avg_disc_unl_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_disc_unl_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_avg_disc_unl_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_l_inst_l_count_order_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_count_order_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_count_order_dvalid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_count_order_last : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_count_order : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummaryWriter_l_inst_l_count_order_bus_wreq_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_count_order_bus_wreq_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_count_order_bus_wreq_addr : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_count_order_bus_wreq_len : STD_LOGIC_VECTOR(BUS_LEN_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_count_order_bus_wdat_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_count_order_bus_wdat_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_count_order_bus_wdat_data : STD_LOGIC_VECTOR(BUS_DATA_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_count_order_bus_wdat_strobe : STD_LOGIC_VECTOR(BUS_DATA_WIDTH/8 - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_count_order_bus_wdat_last : STD_LOGIC;

  SIGNAL PriceSummaryWriter_l_inst_l_count_order_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_count_order_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_count_order_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_count_order_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_count_order_cmd_ctrl : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummaryWriter_l_inst_l_count_order_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummaryWriter_l_inst_l_count_order_unl_valid : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_count_order_unl_ready : STD_LOGIC;
  SIGNAL PriceSummaryWriter_l_inst_l_count_order_unl_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummary_Nucleus_inst_mmio_awvalid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_mmio_awready : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_mmio_awaddr : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummary_Nucleus_inst_mmio_wvalid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_mmio_wready : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_mmio_wdata : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummary_Nucleus_inst_mmio_wstrb : STD_LOGIC_VECTOR(3 DOWNTO 0);
  SIGNAL PriceSummary_Nucleus_inst_mmio_bvalid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_mmio_bready : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_mmio_bresp : STD_LOGIC_VECTOR(1 DOWNTO 0);
  SIGNAL PriceSummary_Nucleus_inst_mmio_arvalid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_mmio_arready : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_mmio_araddr : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummary_Nucleus_inst_mmio_rvalid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_mmio_rready : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_mmio_rdata : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummary_Nucleus_inst_mmio_rresp : STD_LOGIC_VECTOR(1 DOWNTO 0);

  SIGNAL PriceSummary_Nucleus_inst_l_quantity_valid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_quantity_ready : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_quantity_dvalid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_quantity_last : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_quantity : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummary_Nucleus_inst_l_extendedprice_valid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_extendedprice_ready : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_extendedprice_dvalid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_extendedprice_last : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_extendedprice : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummary_Nucleus_inst_l_discount_valid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_discount_ready : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_discount_dvalid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_discount_last : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_discount : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummary_Nucleus_inst_l_tax_valid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_tax_ready : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_tax_dvalid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_tax_last : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_tax : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummary_Nucleus_inst_l_returnflag_valid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_returnflag_ready : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_returnflag_dvalid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_returnflag_last : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_returnflag_length : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummary_Nucleus_inst_l_returnflag_count : STD_LOGIC_VECTOR(0 DOWNTO 0);
  SIGNAL PriceSummary_Nucleus_inst_l_returnflag_chars_valid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_returnflag_chars_ready : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_returnflag_chars_dvalid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_returnflag_chars_last : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_returnflag_chars : STD_LOGIC_VECTOR(7 DOWNTO 0);
  SIGNAL PriceSummary_Nucleus_inst_l_returnflag_chars_count : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummary_Nucleus_inst_l_linestatus_valid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_linestatus_ready : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_linestatus_dvalid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_linestatus_last : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_linestatus_length : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummary_Nucleus_inst_l_linestatus_count : STD_LOGIC_VECTOR(0 DOWNTO 0);
  SIGNAL PriceSummary_Nucleus_inst_l_linestatus_chars_valid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_linestatus_chars_ready : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_linestatus_chars_dvalid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_linestatus_chars_last : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_linestatus_chars : STD_LOGIC_VECTOR(7 DOWNTO 0);
  SIGNAL PriceSummary_Nucleus_inst_l_linestatus_chars_count : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummary_Nucleus_inst_l_shipdate_valid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_shipdate_ready : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_shipdate_dvalid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_shipdate_last : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_shipdate : STD_LOGIC_VECTOR(31 DOWNTO 0);

  SIGNAL PriceSummary_Nucleus_inst_l_quantity_unl_valid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_quantity_unl_ready : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_quantity_unl_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummary_Nucleus_inst_l_extendedprice_unl_valid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_extendedprice_unl_ready : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_extendedprice_unl_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummary_Nucleus_inst_l_discount_unl_valid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_discount_unl_ready : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_discount_unl_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummary_Nucleus_inst_l_tax_unl_valid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_tax_unl_ready : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_tax_unl_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummary_Nucleus_inst_l_returnflag_unl_valid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_returnflag_unl_ready : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_returnflag_unl_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummary_Nucleus_inst_l_linestatus_unl_valid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_linestatus_unl_ready : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_linestatus_unl_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummary_Nucleus_inst_l_shipdate_unl_valid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_shipdate_unl_ready : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_shipdate_unl_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummary_Nucleus_inst_l_quantity_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_quantity_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_quantity_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_Nucleus_inst_l_quantity_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_Nucleus_inst_l_quantity_cmd_ctrl : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_Nucleus_inst_l_quantity_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummary_Nucleus_inst_l_extendedprice_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_extendedprice_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_extendedprice_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_Nucleus_inst_l_extendedprice_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_Nucleus_inst_l_extendedprice_cmd_ctrl : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_Nucleus_inst_l_extendedprice_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummary_Nucleus_inst_l_discount_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_discount_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_discount_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_Nucleus_inst_l_discount_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_Nucleus_inst_l_discount_cmd_ctrl : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_Nucleus_inst_l_discount_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummary_Nucleus_inst_l_tax_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_tax_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_tax_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_Nucleus_inst_l_tax_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_Nucleus_inst_l_tax_cmd_ctrl : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_Nucleus_inst_l_tax_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummary_Nucleus_inst_l_returnflag_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_returnflag_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_returnflag_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_Nucleus_inst_l_returnflag_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_Nucleus_inst_l_returnflag_cmd_ctrl : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH * 2 - 1 DOWNTO 0);
  SIGNAL PriceSummary_Nucleus_inst_l_returnflag_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummary_Nucleus_inst_l_linestatus_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_linestatus_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_linestatus_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_Nucleus_inst_l_linestatus_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_Nucleus_inst_l_linestatus_cmd_ctrl : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH * 2 - 1 DOWNTO 0);
  SIGNAL PriceSummary_Nucleus_inst_l_linestatus_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummary_Nucleus_inst_l_shipdate_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_shipdate_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummary_Nucleus_inst_l_shipdate_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_Nucleus_inst_l_shipdate_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_Nucleus_inst_l_shipdate_cmd_ctrl : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_Nucleus_inst_l_shipdate_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummary_l_inst_l_quantity_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_quantity_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_quantity_dvalid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_quantity_last : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_quantity : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummary_l_inst_l_quantity_bus_rreq_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_quantity_bus_rreq_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_quantity_bus_rreq_addr : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_quantity_bus_rreq_len : STD_LOGIC_VECTOR(BUS_LEN_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_quantity_bus_rdat_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_quantity_bus_rdat_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_quantity_bus_rdat_data : STD_LOGIC_VECTOR(BUS_DATA_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_quantity_bus_rdat_last : STD_LOGIC;

  SIGNAL PriceSummary_l_inst_l_quantity_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_quantity_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_quantity_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_quantity_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_quantity_cmd_ctrl : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_quantity_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummary_l_inst_l_quantity_unl_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_quantity_unl_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_quantity_unl_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummary_l_inst_l_extendedprice_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_extendedprice_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_extendedprice_dvalid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_extendedprice_last : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_extendedprice : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummary_l_inst_l_extendedprice_bus_rreq_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_extendedprice_bus_rreq_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_extendedprice_bus_rreq_addr : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_extendedprice_bus_rreq_len : STD_LOGIC_VECTOR(BUS_LEN_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_extendedprice_bus_rdat_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_extendedprice_bus_rdat_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_extendedprice_bus_rdat_data : STD_LOGIC_VECTOR(BUS_DATA_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_extendedprice_bus_rdat_last : STD_LOGIC;

  SIGNAL PriceSummary_l_inst_l_extendedprice_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_extendedprice_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_extendedprice_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_extendedprice_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_extendedprice_cmd_ctrl : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_extendedprice_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummary_l_inst_l_extendedprice_unl_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_extendedprice_unl_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_extendedprice_unl_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummary_l_inst_l_discount_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_discount_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_discount_dvalid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_discount_last : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_discount : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummary_l_inst_l_discount_bus_rreq_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_discount_bus_rreq_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_discount_bus_rreq_addr : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_discount_bus_rreq_len : STD_LOGIC_VECTOR(BUS_LEN_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_discount_bus_rdat_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_discount_bus_rdat_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_discount_bus_rdat_data : STD_LOGIC_VECTOR(BUS_DATA_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_discount_bus_rdat_last : STD_LOGIC;

  SIGNAL PriceSummary_l_inst_l_discount_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_discount_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_discount_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_discount_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_discount_cmd_ctrl : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_discount_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummary_l_inst_l_discount_unl_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_discount_unl_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_discount_unl_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummary_l_inst_l_tax_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_tax_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_tax_dvalid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_tax_last : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_tax : STD_LOGIC_VECTOR(63 DOWNTO 0);

  SIGNAL PriceSummary_l_inst_l_tax_bus_rreq_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_tax_bus_rreq_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_tax_bus_rreq_addr : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_tax_bus_rreq_len : STD_LOGIC_VECTOR(BUS_LEN_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_tax_bus_rdat_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_tax_bus_rdat_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_tax_bus_rdat_data : STD_LOGIC_VECTOR(BUS_DATA_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_tax_bus_rdat_last : STD_LOGIC;

  SIGNAL PriceSummary_l_inst_l_tax_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_tax_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_tax_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_tax_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_tax_cmd_ctrl : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_tax_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummary_l_inst_l_tax_unl_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_tax_unl_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_tax_unl_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummary_l_inst_l_returnflag_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_returnflag_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_returnflag_dvalid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_returnflag_last : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_returnflag_length : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_returnflag_count : STD_LOGIC_VECTOR(0 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_returnflag_chars_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_returnflag_chars_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_returnflag_chars_dvalid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_returnflag_chars_last : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_returnflag_chars : STD_LOGIC_VECTOR(7 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_returnflag_chars_count : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummary_l_inst_l_returnflag_bus_rreq_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_returnflag_bus_rreq_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_returnflag_bus_rreq_addr : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_returnflag_bus_rreq_len : STD_LOGIC_VECTOR(BUS_LEN_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_returnflag_bus_rdat_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_returnflag_bus_rdat_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_returnflag_bus_rdat_data : STD_LOGIC_VECTOR(BUS_DATA_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_returnflag_bus_rdat_last : STD_LOGIC;

  SIGNAL PriceSummary_l_inst_l_returnflag_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_returnflag_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_returnflag_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_returnflag_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_returnflag_cmd_ctrl : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH * 2 - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_returnflag_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummary_l_inst_l_returnflag_unl_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_returnflag_unl_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_returnflag_unl_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummary_l_inst_l_linestatus_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_linestatus_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_linestatus_dvalid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_linestatus_last : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_linestatus_length : STD_LOGIC_VECTOR(31 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_linestatus_count : STD_LOGIC_VECTOR(0 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_linestatus_chars_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_linestatus_chars_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_linestatus_chars_dvalid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_linestatus_chars_last : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_linestatus_chars : STD_LOGIC_VECTOR(7 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_linestatus_chars_count : STD_LOGIC_VECTOR(0 DOWNTO 0);

  SIGNAL PriceSummary_l_inst_l_linestatus_bus_rreq_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_linestatus_bus_rreq_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_linestatus_bus_rreq_addr : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_linestatus_bus_rreq_len : STD_LOGIC_VECTOR(BUS_LEN_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_linestatus_bus_rdat_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_linestatus_bus_rdat_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_linestatus_bus_rdat_data : STD_LOGIC_VECTOR(BUS_DATA_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_linestatus_bus_rdat_last : STD_LOGIC;

  SIGNAL PriceSummary_l_inst_l_linestatus_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_linestatus_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_linestatus_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_linestatus_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_linestatus_cmd_ctrl : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH * 2 - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_linestatus_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummary_l_inst_l_linestatus_unl_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_linestatus_unl_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_linestatus_unl_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummary_l_inst_l_shipdate_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_shipdate_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_shipdate_dvalid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_shipdate_last : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_shipdate : STD_LOGIC_VECTOR(31 DOWNTO 0);

  SIGNAL PriceSummary_l_inst_l_shipdate_bus_rreq_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_shipdate_bus_rreq_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_shipdate_bus_rreq_addr : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_shipdate_bus_rreq_len : STD_LOGIC_VECTOR(BUS_LEN_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_shipdate_bus_rdat_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_shipdate_bus_rdat_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_shipdate_bus_rdat_data : STD_LOGIC_VECTOR(BUS_DATA_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_shipdate_bus_rdat_last : STD_LOGIC;

  SIGNAL PriceSummary_l_inst_l_shipdate_cmd_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_shipdate_cmd_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_shipdate_cmd_firstIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_shipdate_cmd_lastIdx : STD_LOGIC_VECTOR(INDEX_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_shipdate_cmd_ctrl : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL PriceSummary_l_inst_l_shipdate_cmd_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL PriceSummary_l_inst_l_shipdate_unl_valid : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_shipdate_unl_ready : STD_LOGIC;
  SIGNAL PriceSummary_l_inst_l_shipdate_unl_tag : STD_LOGIC_VECTOR(TAG_WIDTH - 1 DOWNTO 0);

  SIGNAL RDAW64DW512LW8BS1BM16_inst_mst_rreq_valid : STD_LOGIC;
  SIGNAL RDAW64DW512LW8BS1BM16_inst_mst_rreq_ready : STD_LOGIC;
  SIGNAL RDAW64DW512LW8BS1BM16_inst_mst_rreq_addr : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL RDAW64DW512LW8BS1BM16_inst_mst_rreq_len : STD_LOGIC_VECTOR(BUS_LEN_WIDTH - 1 DOWNTO 0);
  SIGNAL RDAW64DW512LW8BS1BM16_inst_mst_rdat_valid : STD_LOGIC;
  SIGNAL RDAW64DW512LW8BS1BM16_inst_mst_rdat_ready : STD_LOGIC;
  SIGNAL RDAW64DW512LW8BS1BM16_inst_mst_rdat_data : STD_LOGIC_VECTOR(BUS_DATA_WIDTH - 1 DOWNTO 0);
  SIGNAL RDAW64DW512LW8BS1BM16_inst_mst_rdat_last : STD_LOGIC;

  SIGNAL RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid : STD_LOGIC_VECTOR(6 DOWNTO 0);
  SIGNAL RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready : STD_LOGIC_VECTOR(6 DOWNTO 0);
  SIGNAL RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr : STD_LOGIC_VECTOR(7 * BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len : STD_LOGIC_VECTOR(7 * BUS_LEN_WIDTH - 1 DOWNTO 0);
  SIGNAL RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid : STD_LOGIC_VECTOR(6 DOWNTO 0);
  SIGNAL RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready : STD_LOGIC_VECTOR(6 DOWNTO 0);
  SIGNAL RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data : STD_LOGIC_VECTOR(7 * BUS_DATA_WIDTH - 1 DOWNTO 0);
  SIGNAL RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last : STD_LOGIC_VECTOR(6 DOWNTO 0);

  SIGNAL WRAW64DW512LW8BS1BM16_inst_mst_wreq_valid : STD_LOGIC;
  SIGNAL WRAW64DW512LW8BS1BM16_inst_mst_wreq_ready : STD_LOGIC;
  SIGNAL WRAW64DW512LW8BS1BM16_inst_mst_wreq_addr : STD_LOGIC_VECTOR(BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL WRAW64DW512LW8BS1BM16_inst_mst_wreq_len : STD_LOGIC_VECTOR(BUS_LEN_WIDTH - 1 DOWNTO 0);
  SIGNAL WRAW64DW512LW8BS1BM16_inst_mst_wdat_valid : STD_LOGIC;
  SIGNAL WRAW64DW512LW8BS1BM16_inst_mst_wdat_ready : STD_LOGIC;
  SIGNAL WRAW64DW512LW8BS1BM16_inst_mst_wdat_data : STD_LOGIC_VECTOR(BUS_DATA_WIDTH - 1 DOWNTO 0);
  SIGNAL WRAW64DW512LW8BS1BM16_inst_mst_wdat_strobe : STD_LOGIC_VECTOR(BUS_DATA_WIDTH/8 - 1 DOWNTO 0);
  SIGNAL WRAW64DW512LW8BS1BM16_inst_mst_wdat_last : STD_LOGIC;

  SIGNAL WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid : STD_LOGIC_VECTOR(9 DOWNTO 0);
  SIGNAL WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready : STD_LOGIC_VECTOR(9 DOWNTO 0);
  SIGNAL WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr : STD_LOGIC_VECTOR(10 * BUS_ADDR_WIDTH - 1 DOWNTO 0);
  SIGNAL WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len : STD_LOGIC_VECTOR(10 * BUS_LEN_WIDTH - 1 DOWNTO 0);
  SIGNAL WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid : STD_LOGIC_VECTOR(9 DOWNTO 0);
  SIGNAL WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready : STD_LOGIC_VECTOR(9 DOWNTO 0);
  SIGNAL WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data : STD_LOGIC_VECTOR(10 * BUS_DATA_WIDTH - 1 DOWNTO 0);
  SIGNAL WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe : STD_LOGIC_VECTOR(10 * BUS_DATA_WIDTH/8 - 1 DOWNTO 0);
  SIGNAL WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last : STD_LOGIC_VECTOR(9 DOWNTO 0);
BEGIN
  PriceSummary_Nucleus_inst : PriceSummary_Nucleus
  GENERIC MAP(
    INDEX_WIDTH => INDEX_WIDTH,
    TAG_WIDTH => TAG_WIDTH,
    L_QUANTITY_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_EXTENDEDPRICE_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_DISCOUNT_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_TAX_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_RETURNFLAG_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_LINESTATUS_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_SHIPDATE_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_RETURNFLAG_O_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_LINESTATUS_O_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_SUM_QTY_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_SUM_BASE_PRICE_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_SUM_DISC_PRICE_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_SUM_CHARGE_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_AVG_QTY_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_AVG_PRICE_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_AVG_DISC_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_COUNT_ORDER_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH
  )
  PORT MAP(
    kcd_clk => kcd_clk,
    kcd_reset => kcd_reset,
    mmio_awvalid => PriceSummary_Nucleus_inst_mmio_awvalid,
    mmio_awready => PriceSummary_Nucleus_inst_mmio_awready,
    mmio_awaddr => PriceSummary_Nucleus_inst_mmio_awaddr,
    mmio_wvalid => PriceSummary_Nucleus_inst_mmio_wvalid,
    mmio_wready => PriceSummary_Nucleus_inst_mmio_wready,
    mmio_wdata => PriceSummary_Nucleus_inst_mmio_wdata,
    mmio_wstrb => PriceSummary_Nucleus_inst_mmio_wstrb,
    mmio_bvalid => PriceSummary_Nucleus_inst_mmio_bvalid,
    mmio_bready => PriceSummary_Nucleus_inst_mmio_bready,
    mmio_bresp => PriceSummary_Nucleus_inst_mmio_bresp,
    mmio_arvalid => PriceSummary_Nucleus_inst_mmio_arvalid,
    mmio_arready => PriceSummary_Nucleus_inst_mmio_arready,
    mmio_araddr => PriceSummary_Nucleus_inst_mmio_araddr,
    mmio_rvalid => PriceSummary_Nucleus_inst_mmio_rvalid,
    mmio_rready => PriceSummary_Nucleus_inst_mmio_rready,
    mmio_rdata => PriceSummary_Nucleus_inst_mmio_rdata,
    mmio_rresp => PriceSummary_Nucleus_inst_mmio_rresp,
    l_quantity_valid => PriceSummary_Nucleus_inst_l_quantity_valid,
    l_quantity_ready => PriceSummary_Nucleus_inst_l_quantity_ready,
    l_quantity_dvalid => PriceSummary_Nucleus_inst_l_quantity_dvalid,
    l_quantity_last => PriceSummary_Nucleus_inst_l_quantity_last,
    l_quantity => PriceSummary_Nucleus_inst_l_quantity,
    l_extendedprice_valid => PriceSummary_Nucleus_inst_l_extendedprice_valid,
    l_extendedprice_ready => PriceSummary_Nucleus_inst_l_extendedprice_ready,
    l_extendedprice_dvalid => PriceSummary_Nucleus_inst_l_extendedprice_dvalid,
    l_extendedprice_last => PriceSummary_Nucleus_inst_l_extendedprice_last,
    l_extendedprice => PriceSummary_Nucleus_inst_l_extendedprice,
    l_discount_valid => PriceSummary_Nucleus_inst_l_discount_valid,
    l_discount_ready => PriceSummary_Nucleus_inst_l_discount_ready,
    l_discount_dvalid => PriceSummary_Nucleus_inst_l_discount_dvalid,
    l_discount_last => PriceSummary_Nucleus_inst_l_discount_last,
    l_discount => PriceSummary_Nucleus_inst_l_discount,
    l_tax_valid => PriceSummary_Nucleus_inst_l_tax_valid,
    l_tax_ready => PriceSummary_Nucleus_inst_l_tax_ready,
    l_tax_dvalid => PriceSummary_Nucleus_inst_l_tax_dvalid,
    l_tax_last => PriceSummary_Nucleus_inst_l_tax_last,
    l_tax => PriceSummary_Nucleus_inst_l_tax,
    l_returnflag_valid => PriceSummary_Nucleus_inst_l_returnflag_valid,
    l_returnflag_ready => PriceSummary_Nucleus_inst_l_returnflag_ready,
    l_returnflag_dvalid => PriceSummary_Nucleus_inst_l_returnflag_dvalid,
    l_returnflag_last => PriceSummary_Nucleus_inst_l_returnflag_last,
    l_returnflag_length => PriceSummary_Nucleus_inst_l_returnflag_length,
    l_returnflag_count => PriceSummary_Nucleus_inst_l_returnflag_count,
    l_returnflag_chars_valid => PriceSummary_Nucleus_inst_l_returnflag_chars_valid,
    l_returnflag_chars_ready => PriceSummary_Nucleus_inst_l_returnflag_chars_ready,
    l_returnflag_chars_dvalid => PriceSummary_Nucleus_inst_l_returnflag_chars_dvalid,
    l_returnflag_chars_last => PriceSummary_Nucleus_inst_l_returnflag_chars_last,
    l_returnflag_chars => PriceSummary_Nucleus_inst_l_returnflag_chars,
    l_returnflag_chars_count => PriceSummary_Nucleus_inst_l_returnflag_chars_count,
    l_linestatus_valid => PriceSummary_Nucleus_inst_l_linestatus_valid,
    l_linestatus_ready => PriceSummary_Nucleus_inst_l_linestatus_ready,
    l_linestatus_dvalid => PriceSummary_Nucleus_inst_l_linestatus_dvalid,
    l_linestatus_last => PriceSummary_Nucleus_inst_l_linestatus_last,
    l_linestatus_length => PriceSummary_Nucleus_inst_l_linestatus_length,
    l_linestatus_count => PriceSummary_Nucleus_inst_l_linestatus_count,
    l_linestatus_chars_valid => PriceSummary_Nucleus_inst_l_linestatus_chars_valid,
    l_linestatus_chars_ready => PriceSummary_Nucleus_inst_l_linestatus_chars_ready,
    l_linestatus_chars_dvalid => PriceSummary_Nucleus_inst_l_linestatus_chars_dvalid,
    l_linestatus_chars_last => PriceSummary_Nucleus_inst_l_linestatus_chars_last,
    l_linestatus_chars => PriceSummary_Nucleus_inst_l_linestatus_chars,
    l_linestatus_chars_count => PriceSummary_Nucleus_inst_l_linestatus_chars_count,
    l_shipdate_valid => PriceSummary_Nucleus_inst_l_shipdate_valid,
    l_shipdate_ready => PriceSummary_Nucleus_inst_l_shipdate_ready,
    l_shipdate_dvalid => PriceSummary_Nucleus_inst_l_shipdate_dvalid,
    l_shipdate_last => PriceSummary_Nucleus_inst_l_shipdate_last,
    l_shipdate => PriceSummary_Nucleus_inst_l_shipdate,
    l_quantity_unl_valid => PriceSummary_Nucleus_inst_l_quantity_unl_valid,
    l_quantity_unl_ready => PriceSummary_Nucleus_inst_l_quantity_unl_ready,
    l_quantity_unl_tag => PriceSummary_Nucleus_inst_l_quantity_unl_tag,
    l_extendedprice_unl_valid => PriceSummary_Nucleus_inst_l_extendedprice_unl_valid,
    l_extendedprice_unl_ready => PriceSummary_Nucleus_inst_l_extendedprice_unl_ready,
    l_extendedprice_unl_tag => PriceSummary_Nucleus_inst_l_extendedprice_unl_tag,
    l_discount_unl_valid => PriceSummary_Nucleus_inst_l_discount_unl_valid,
    l_discount_unl_ready => PriceSummary_Nucleus_inst_l_discount_unl_ready,
    l_discount_unl_tag => PriceSummary_Nucleus_inst_l_discount_unl_tag,
    l_tax_unl_valid => PriceSummary_Nucleus_inst_l_tax_unl_valid,
    l_tax_unl_ready => PriceSummary_Nucleus_inst_l_tax_unl_ready,
    l_tax_unl_tag => PriceSummary_Nucleus_inst_l_tax_unl_tag,
    l_returnflag_unl_valid => PriceSummary_Nucleus_inst_l_returnflag_unl_valid,
    l_returnflag_unl_ready => PriceSummary_Nucleus_inst_l_returnflag_unl_ready,
    l_returnflag_unl_tag => PriceSummary_Nucleus_inst_l_returnflag_unl_tag,
    l_linestatus_unl_valid => PriceSummary_Nucleus_inst_l_linestatus_unl_valid,
    l_linestatus_unl_ready => PriceSummary_Nucleus_inst_l_linestatus_unl_ready,
    l_linestatus_unl_tag => PriceSummary_Nucleus_inst_l_linestatus_unl_tag,
    l_shipdate_unl_valid => PriceSummary_Nucleus_inst_l_shipdate_unl_valid,
    l_shipdate_unl_ready => PriceSummary_Nucleus_inst_l_shipdate_unl_ready,
    l_shipdate_unl_tag => PriceSummary_Nucleus_inst_l_shipdate_unl_tag,
    l_quantity_cmd_valid => PriceSummary_Nucleus_inst_l_quantity_cmd_valid,
    l_quantity_cmd_ready => PriceSummary_Nucleus_inst_l_quantity_cmd_ready,
    l_quantity_cmd_firstIdx => PriceSummary_Nucleus_inst_l_quantity_cmd_firstIdx,
    l_quantity_cmd_lastIdx => PriceSummary_Nucleus_inst_l_quantity_cmd_lastIdx,
    l_quantity_cmd_ctrl => PriceSummary_Nucleus_inst_l_quantity_cmd_ctrl,
    l_quantity_cmd_tag => PriceSummary_Nucleus_inst_l_quantity_cmd_tag,
    l_extendedprice_cmd_valid => PriceSummary_Nucleus_inst_l_extendedprice_cmd_valid,
    l_extendedprice_cmd_ready => PriceSummary_Nucleus_inst_l_extendedprice_cmd_ready,
    l_extendedprice_cmd_firstIdx => PriceSummary_Nucleus_inst_l_extendedprice_cmd_firstIdx,
    l_extendedprice_cmd_lastIdx => PriceSummary_Nucleus_inst_l_extendedprice_cmd_lastIdx,
    l_extendedprice_cmd_ctrl => PriceSummary_Nucleus_inst_l_extendedprice_cmd_ctrl,
    l_extendedprice_cmd_tag => PriceSummary_Nucleus_inst_l_extendedprice_cmd_tag,
    l_discount_cmd_valid => PriceSummary_Nucleus_inst_l_discount_cmd_valid,
    l_discount_cmd_ready => PriceSummary_Nucleus_inst_l_discount_cmd_ready,
    l_discount_cmd_firstIdx => PriceSummary_Nucleus_inst_l_discount_cmd_firstIdx,
    l_discount_cmd_lastIdx => PriceSummary_Nucleus_inst_l_discount_cmd_lastIdx,
    l_discount_cmd_ctrl => PriceSummary_Nucleus_inst_l_discount_cmd_ctrl,
    l_discount_cmd_tag => PriceSummary_Nucleus_inst_l_discount_cmd_tag,
    l_tax_cmd_valid => PriceSummary_Nucleus_inst_l_tax_cmd_valid,
    l_tax_cmd_ready => PriceSummary_Nucleus_inst_l_tax_cmd_ready,
    l_tax_cmd_firstIdx => PriceSummary_Nucleus_inst_l_tax_cmd_firstIdx,
    l_tax_cmd_lastIdx => PriceSummary_Nucleus_inst_l_tax_cmd_lastIdx,
    l_tax_cmd_ctrl => PriceSummary_Nucleus_inst_l_tax_cmd_ctrl,
    l_tax_cmd_tag => PriceSummary_Nucleus_inst_l_tax_cmd_tag,
    l_returnflag_cmd_valid => PriceSummary_Nucleus_inst_l_returnflag_cmd_valid,
    l_returnflag_cmd_ready => PriceSummary_Nucleus_inst_l_returnflag_cmd_ready,
    l_returnflag_cmd_firstIdx => PriceSummary_Nucleus_inst_l_returnflag_cmd_firstIdx,
    l_returnflag_cmd_lastIdx => PriceSummary_Nucleus_inst_l_returnflag_cmd_lastIdx,
    l_returnflag_cmd_ctrl => PriceSummary_Nucleus_inst_l_returnflag_cmd_ctrl,
    l_returnflag_cmd_tag => PriceSummary_Nucleus_inst_l_returnflag_cmd_tag,
    l_linestatus_cmd_valid => PriceSummary_Nucleus_inst_l_linestatus_cmd_valid,
    l_linestatus_cmd_ready => PriceSummary_Nucleus_inst_l_linestatus_cmd_ready,
    l_linestatus_cmd_firstIdx => PriceSummary_Nucleus_inst_l_linestatus_cmd_firstIdx,
    l_linestatus_cmd_lastIdx => PriceSummary_Nucleus_inst_l_linestatus_cmd_lastIdx,
    l_linestatus_cmd_ctrl => PriceSummary_Nucleus_inst_l_linestatus_cmd_ctrl,
    l_linestatus_cmd_tag => PriceSummary_Nucleus_inst_l_linestatus_cmd_tag,
    l_shipdate_cmd_valid => PriceSummary_Nucleus_inst_l_shipdate_cmd_valid,
    l_shipdate_cmd_ready => PriceSummary_Nucleus_inst_l_shipdate_cmd_ready,
    l_shipdate_cmd_firstIdx => PriceSummary_Nucleus_inst_l_shipdate_cmd_firstIdx,
    l_shipdate_cmd_lastIdx => PriceSummary_Nucleus_inst_l_shipdate_cmd_lastIdx,
    l_shipdate_cmd_ctrl => PriceSummary_Nucleus_inst_l_shipdate_cmd_ctrl,
    l_shipdate_cmd_tag => PriceSummary_Nucleus_inst_l_shipdate_cmd_tag,
    l_returnflag_o_valid => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_valid,
    l_returnflag_o_ready => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_ready,
    l_returnflag_o_dvalid => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_dvalid,
    l_returnflag_o_last => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_last,
    l_returnflag_o_length => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_length,
    l_returnflag_o_count => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_count,
    l_returnflag_o_chars_valid => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_valid,
    l_returnflag_o_chars_ready => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_ready,
    l_returnflag_o_chars_dvalid => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_dvalid,
    l_returnflag_o_chars_last => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_last,
    l_returnflag_o_chars => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars,
    l_returnflag_o_chars_count => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_count,
    l_linestatus_o_valid => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_valid,
    l_linestatus_o_ready => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_ready,
    l_linestatus_o_dvalid => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_dvalid,
    l_linestatus_o_last => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_last,
    l_linestatus_o_length => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_length,
    l_linestatus_o_count => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_count,
    l_linestatus_o_chars_valid => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_valid,
    l_linestatus_o_chars_ready => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_ready,
    l_linestatus_o_chars_dvalid => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_dvalid,
    l_linestatus_o_chars_last => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_last,
    l_linestatus_o_chars => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars,
    l_linestatus_o_chars_count => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_count,
    l_sum_qty_valid => PriceSummaryWriter_Nucleus_inst_l_sum_qty_valid,
    l_sum_qty_ready => PriceSummaryWriter_Nucleus_inst_l_sum_qty_ready,
    l_sum_qty_dvalid => PriceSummaryWriter_Nucleus_inst_l_sum_qty_dvalid,
    l_sum_qty_last => PriceSummaryWriter_Nucleus_inst_l_sum_qty_last,
    l_sum_qty => PriceSummaryWriter_Nucleus_inst_l_sum_qty,
    l_sum_base_price_valid => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_valid,
    l_sum_base_price_ready => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_ready,
    l_sum_base_price_dvalid => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_dvalid,
    l_sum_base_price_last => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_last,
    l_sum_base_price => PriceSummaryWriter_Nucleus_inst_l_sum_base_price,
    l_sum_disc_price_valid => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_valid,
    l_sum_disc_price_ready => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_ready,
    l_sum_disc_price_dvalid => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_dvalid,
    l_sum_disc_price_last => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_last,
    l_sum_disc_price => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price,
    l_sum_charge_valid => PriceSummaryWriter_Nucleus_inst_l_sum_charge_valid,
    l_sum_charge_ready => PriceSummaryWriter_Nucleus_inst_l_sum_charge_ready,
    l_sum_charge_dvalid => PriceSummaryWriter_Nucleus_inst_l_sum_charge_dvalid,
    l_sum_charge_last => PriceSummaryWriter_Nucleus_inst_l_sum_charge_last,
    l_sum_charge => PriceSummaryWriter_Nucleus_inst_l_sum_charge,
    l_avg_qty_valid => PriceSummaryWriter_Nucleus_inst_l_avg_qty_valid,
    l_avg_qty_ready => PriceSummaryWriter_Nucleus_inst_l_avg_qty_ready,
    l_avg_qty_dvalid => PriceSummaryWriter_Nucleus_inst_l_avg_qty_dvalid,
    l_avg_qty_last => PriceSummaryWriter_Nucleus_inst_l_avg_qty_last,
    l_avg_qty => PriceSummaryWriter_Nucleus_inst_l_avg_qty,
    l_avg_price_valid => PriceSummaryWriter_Nucleus_inst_l_avg_price_valid,
    l_avg_price_ready => PriceSummaryWriter_Nucleus_inst_l_avg_price_ready,
    l_avg_price_dvalid => PriceSummaryWriter_Nucleus_inst_l_avg_price_dvalid,
    l_avg_price_last => PriceSummaryWriter_Nucleus_inst_l_avg_price_last,
    l_avg_price => PriceSummaryWriter_Nucleus_inst_l_avg_price,
    l_avg_disc_valid => PriceSummaryWriter_Nucleus_inst_l_avg_disc_valid,
    l_avg_disc_ready => PriceSummaryWriter_Nucleus_inst_l_avg_disc_ready,
    l_avg_disc_dvalid => PriceSummaryWriter_Nucleus_inst_l_avg_disc_dvalid,
    l_avg_disc_last => PriceSummaryWriter_Nucleus_inst_l_avg_disc_last,
    l_avg_disc => PriceSummaryWriter_Nucleus_inst_l_avg_disc,
    l_count_order_valid => PriceSummaryWriter_Nucleus_inst_l_count_order_valid,
    l_count_order_ready => PriceSummaryWriter_Nucleus_inst_l_count_order_ready,
    l_count_order_dvalid => PriceSummaryWriter_Nucleus_inst_l_count_order_dvalid,
    l_count_order_last => PriceSummaryWriter_Nucleus_inst_l_count_order_last,
    l_count_order => PriceSummaryWriter_Nucleus_inst_l_count_order,
    l_returnflag_o_unl_valid => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_unl_valid,
    l_returnflag_o_unl_ready => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_unl_ready,
    l_returnflag_o_unl_tag => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_unl_tag,
    l_linestatus_o_unl_valid => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_unl_valid,
    l_linestatus_o_unl_ready => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_unl_ready,
    l_linestatus_o_unl_tag => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_unl_tag,
    l_sum_qty_unl_valid => PriceSummaryWriter_Nucleus_inst_l_sum_qty_unl_valid,
    l_sum_qty_unl_ready => PriceSummaryWriter_Nucleus_inst_l_sum_qty_unl_ready,
    l_sum_qty_unl_tag => PriceSummaryWriter_Nucleus_inst_l_sum_qty_unl_tag,
    l_sum_base_price_unl_valid => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_unl_valid,
    l_sum_base_price_unl_ready => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_unl_ready,
    l_sum_base_price_unl_tag => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_unl_tag,
    l_sum_disc_price_unl_valid => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_unl_valid,
    l_sum_disc_price_unl_ready => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_unl_ready,
    l_sum_disc_price_unl_tag => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_unl_tag,
    l_sum_charge_unl_valid => PriceSummaryWriter_Nucleus_inst_l_sum_charge_unl_valid,
    l_sum_charge_unl_ready => PriceSummaryWriter_Nucleus_inst_l_sum_charge_unl_ready,
    l_sum_charge_unl_tag => PriceSummaryWriter_Nucleus_inst_l_sum_charge_unl_tag,
    l_avg_qty_unl_valid => PriceSummaryWriter_Nucleus_inst_l_avg_qty_unl_valid,
    l_avg_qty_unl_ready => PriceSummaryWriter_Nucleus_inst_l_avg_qty_unl_ready,
    l_avg_qty_unl_tag => PriceSummaryWriter_Nucleus_inst_l_avg_qty_unl_tag,
    l_avg_price_unl_valid => PriceSummaryWriter_Nucleus_inst_l_avg_price_unl_valid,
    l_avg_price_unl_ready => PriceSummaryWriter_Nucleus_inst_l_avg_price_unl_ready,
    l_avg_price_unl_tag => PriceSummaryWriter_Nucleus_inst_l_avg_price_unl_tag,
    l_avg_disc_unl_valid => PriceSummaryWriter_Nucleus_inst_l_avg_disc_unl_valid,
    l_avg_disc_unl_ready => PriceSummaryWriter_Nucleus_inst_l_avg_disc_unl_ready,
    l_avg_disc_unl_tag => PriceSummaryWriter_Nucleus_inst_l_avg_disc_unl_tag,
    l_count_order_unl_valid => PriceSummaryWriter_Nucleus_inst_l_count_order_unl_valid,
    l_count_order_unl_ready => PriceSummaryWriter_Nucleus_inst_l_count_order_unl_ready,
    l_count_order_unl_tag => PriceSummaryWriter_Nucleus_inst_l_count_order_unl_tag,
    l_returnflag_o_cmd_valid => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_valid,
    l_returnflag_o_cmd_ready => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_ready,
    l_returnflag_o_cmd_firstIdx => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_firstIdx,
    l_returnflag_o_cmd_lastIdx => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_lastIdx,
    l_returnflag_o_cmd_ctrl => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_ctrl,
    l_returnflag_o_cmd_tag => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_tag,
    l_linestatus_o_cmd_valid => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_valid,
    l_linestatus_o_cmd_ready => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_ready,
    l_linestatus_o_cmd_firstIdx => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_firstIdx,
    l_linestatus_o_cmd_lastIdx => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_lastIdx,
    l_linestatus_o_cmd_ctrl => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_ctrl,
    l_linestatus_o_cmd_tag => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_tag,
    l_sum_qty_cmd_valid => PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_valid,
    l_sum_qty_cmd_ready => PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_ready,
    l_sum_qty_cmd_firstIdx => PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_firstIdx,
    l_sum_qty_cmd_lastIdx => PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_lastIdx,
    l_sum_qty_cmd_ctrl => PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_ctrl,
    l_sum_qty_cmd_tag => PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_tag,
    l_sum_base_price_cmd_valid => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_valid,
    l_sum_base_price_cmd_ready => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_ready,
    l_sum_base_price_cmd_firstIdx => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_firstIdx,
    l_sum_base_price_cmd_lastIdx => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_lastIdx,
    l_sum_base_price_cmd_ctrl => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_ctrl,
    l_sum_base_price_cmd_tag => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_tag,
    l_sum_disc_price_cmd_valid => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_valid,
    l_sum_disc_price_cmd_ready => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_ready,
    l_sum_disc_price_cmd_firstIdx => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_firstIdx,
    l_sum_disc_price_cmd_lastIdx => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_lastIdx,
    l_sum_disc_price_cmd_ctrl => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_ctrl,
    l_sum_disc_price_cmd_tag => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_tag,
    l_sum_charge_cmd_valid => PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_valid,
    l_sum_charge_cmd_ready => PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_ready,
    l_sum_charge_cmd_firstIdx => PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_firstIdx,
    l_sum_charge_cmd_lastIdx => PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_lastIdx,
    l_sum_charge_cmd_ctrl => PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_ctrl,
    l_sum_charge_cmd_tag => PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_tag,
    l_avg_qty_cmd_valid => PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_valid,
    l_avg_qty_cmd_ready => PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_ready,
    l_avg_qty_cmd_firstIdx => PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_firstIdx,
    l_avg_qty_cmd_lastIdx => PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_lastIdx,
    l_avg_qty_cmd_ctrl => PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_ctrl,
    l_avg_qty_cmd_tag => PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_tag,
    l_avg_price_cmd_valid => PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_valid,
    l_avg_price_cmd_ready => PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_ready,
    l_avg_price_cmd_firstIdx => PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_firstIdx,
    l_avg_price_cmd_lastIdx => PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_lastIdx,
    l_avg_price_cmd_ctrl => PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_ctrl,
    l_avg_price_cmd_tag => PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_tag,
    l_avg_disc_cmd_valid => PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_valid,
    l_avg_disc_cmd_ready => PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_ready,
    l_avg_disc_cmd_firstIdx => PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_firstIdx,
    l_avg_disc_cmd_lastIdx => PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_lastIdx,
    l_avg_disc_cmd_ctrl => PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_ctrl,
    l_avg_disc_cmd_tag => PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_tag,
    l_count_order_cmd_valid => PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_valid,
    l_count_order_cmd_ready => PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_ready,
    l_count_order_cmd_firstIdx => PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_firstIdx,
    l_count_order_cmd_lastIdx => PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_lastIdx,
    l_count_order_cmd_ctrl => PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_ctrl,
    l_count_order_cmd_tag => PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_tag
  );

  PriceSummary_l_inst : PriceSummary_l
  GENERIC MAP(
    INDEX_WIDTH => INDEX_WIDTH,
    TAG_WIDTH => TAG_WIDTH,
    L_QUANTITY_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_QUANTITY_BUS_DATA_WIDTH => BUS_DATA_WIDTH,
    L_QUANTITY_BUS_LEN_WIDTH => BUS_LEN_WIDTH,
    L_QUANTITY_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
    L_QUANTITY_BUS_BURST_MAX_LEN => BUS_BURST_MAX_LEN,
    L_EXTENDEDPRICE_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_EXTENDEDPRICE_BUS_DATA_WIDTH => BUS_DATA_WIDTH,
    L_EXTENDEDPRICE_BUS_LEN_WIDTH => BUS_LEN_WIDTH,
    L_EXTENDEDPRICE_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
    L_EXTENDEDPRICE_BUS_BURST_MAX_LEN => BUS_BURST_MAX_LEN,
    L_DISCOUNT_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_DISCOUNT_BUS_DATA_WIDTH => BUS_DATA_WIDTH,
    L_DISCOUNT_BUS_LEN_WIDTH => BUS_LEN_WIDTH,
    L_DISCOUNT_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
    L_DISCOUNT_BUS_BURST_MAX_LEN => BUS_BURST_MAX_LEN,
    L_TAX_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_TAX_BUS_DATA_WIDTH => BUS_DATA_WIDTH,
    L_TAX_BUS_LEN_WIDTH => BUS_LEN_WIDTH,
    L_TAX_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
    L_TAX_BUS_BURST_MAX_LEN => BUS_BURST_MAX_LEN,
    L_RETURNFLAG_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_RETURNFLAG_BUS_DATA_WIDTH => BUS_DATA_WIDTH,
    L_RETURNFLAG_BUS_LEN_WIDTH => BUS_LEN_WIDTH,
    L_RETURNFLAG_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
    L_RETURNFLAG_BUS_BURST_MAX_LEN => BUS_BURST_MAX_LEN,
    L_LINESTATUS_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_LINESTATUS_BUS_DATA_WIDTH => BUS_DATA_WIDTH,
    L_LINESTATUS_BUS_LEN_WIDTH => BUS_LEN_WIDTH,
    L_LINESTATUS_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
    L_LINESTATUS_BUS_BURST_MAX_LEN => BUS_BURST_MAX_LEN,
    L_SHIPDATE_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_SHIPDATE_BUS_DATA_WIDTH => BUS_DATA_WIDTH,
    L_SHIPDATE_BUS_LEN_WIDTH => BUS_LEN_WIDTH,
    L_SHIPDATE_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
    L_SHIPDATE_BUS_BURST_MAX_LEN => BUS_BURST_MAX_LEN,
    L_RETURNFLAG_O_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_RETURNFLAG_O_BUS_DATA_WIDTH => BUS_DATA_WIDTH,
    L_RETURNFLAG_O_BUS_LEN_WIDTH => BUS_LEN_WIDTH,
    L_RETURNFLAG_O_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
    L_RETURNFLAG_O_BUS_BURST_MAX_LEN => BUS_BURST_MAX_LEN,
    L_LINESTATUS_O_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_LINESTATUS_O_BUS_DATA_WIDTH => BUS_DATA_WIDTH,
    L_LINESTATUS_O_BUS_LEN_WIDTH => BUS_LEN_WIDTH,
    L_LINESTATUS_O_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
    L_LINESTATUS_O_BUS_BURST_MAX_LEN => BUS_BURST_MAX_LEN,
    L_SUM_QTY_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_SUM_QTY_BUS_DATA_WIDTH => BUS_DATA_WIDTH,
    L_SUM_QTY_BUS_LEN_WIDTH => BUS_LEN_WIDTH,
    L_SUM_QTY_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
    L_SUM_QTY_BUS_BURST_MAX_LEN => BUS_BURST_MAX_LEN,
    L_SUM_BASE_PRICE_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_SUM_BASE_PRICE_BUS_DATA_WIDTH => BUS_DATA_WIDTH,
    L_SUM_BASE_PRICE_BUS_LEN_WIDTH => BUS_LEN_WIDTH,
    L_SUM_BASE_PRICE_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
    L_SUM_BASE_PRICE_BUS_BURST_MAX_LEN => BUS_BURST_MAX_LEN,
    L_SUM_DISC_PRICE_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_SUM_DISC_PRICE_BUS_DATA_WIDTH => BUS_DATA_WIDTH,
    L_SUM_DISC_PRICE_BUS_LEN_WIDTH => BUS_LEN_WIDTH,
    L_SUM_DISC_PRICE_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
    L_SUM_DISC_PRICE_BUS_BURST_MAX_LEN => BUS_BURST_MAX_LEN,
    L_SUM_CHARGE_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_SUM_CHARGE_BUS_DATA_WIDTH => BUS_DATA_WIDTH,
    L_SUM_CHARGE_BUS_LEN_WIDTH => BUS_LEN_WIDTH,
    L_SUM_CHARGE_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
    L_SUM_CHARGE_BUS_BURST_MAX_LEN => BUS_BURST_MAX_LEN,
    L_AVG_QTY_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_AVG_QTY_BUS_DATA_WIDTH => BUS_DATA_WIDTH,
    L_AVG_QTY_BUS_LEN_WIDTH => BUS_LEN_WIDTH,
    L_AVG_QTY_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
    L_AVG_QTY_BUS_BURST_MAX_LEN => BUS_BURST_MAX_LEN,
    L_AVG_PRICE_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_AVG_PRICE_BUS_DATA_WIDTH => BUS_DATA_WIDTH,
    L_AVG_PRICE_BUS_LEN_WIDTH => BUS_LEN_WIDTH,
    L_AVG_PRICE_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
    L_AVG_PRICE_BUS_BURST_MAX_LEN => BUS_BURST_MAX_LEN,
    L_AVG_DISC_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_AVG_DISC_BUS_DATA_WIDTH => BUS_DATA_WIDTH,
    L_AVG_DISC_BUS_LEN_WIDTH => BUS_LEN_WIDTH,
    L_AVG_DISC_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
    L_AVG_DISC_BUS_BURST_MAX_LEN => BUS_BURST_MAX_LEN,
    L_COUNT_ORDER_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    L_COUNT_ORDER_BUS_DATA_WIDTH => BUS_DATA_WIDTH,
    L_COUNT_ORDER_BUS_LEN_WIDTH => BUS_LEN_WIDTH,
    L_COUNT_ORDER_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
    L_COUNT_ORDER_BUS_BURST_MAX_LEN => BUS_BURST_MAX_LEN
  )
  PORT MAP(
    bcd_clk => bcd_clk,
    bcd_reset => bcd_reset,
    kcd_clk => kcd_clk,
    kcd_reset => kcd_reset,
    l_quantity_valid => PriceSummary_l_inst_l_quantity_valid,
    l_quantity_ready => PriceSummary_l_inst_l_quantity_ready,
    l_quantity_dvalid => PriceSummary_l_inst_l_quantity_dvalid,
    l_quantity_last => PriceSummary_l_inst_l_quantity_last,
    l_quantity => PriceSummary_l_inst_l_quantity,
    l_quantity_bus_rreq_valid => PriceSummary_l_inst_l_quantity_bus_rreq_valid,
    l_quantity_bus_rreq_ready => PriceSummary_l_inst_l_quantity_bus_rreq_ready,
    l_quantity_bus_rreq_addr => PriceSummary_l_inst_l_quantity_bus_rreq_addr,
    l_quantity_bus_rreq_len => PriceSummary_l_inst_l_quantity_bus_rreq_len,
    l_quantity_bus_rdat_valid => PriceSummary_l_inst_l_quantity_bus_rdat_valid,
    l_quantity_bus_rdat_ready => PriceSummary_l_inst_l_quantity_bus_rdat_ready,
    l_quantity_bus_rdat_data => PriceSummary_l_inst_l_quantity_bus_rdat_data,
    l_quantity_bus_rdat_last => PriceSummary_l_inst_l_quantity_bus_rdat_last,
    l_quantity_cmd_valid => PriceSummary_l_inst_l_quantity_cmd_valid,
    l_quantity_cmd_ready => PriceSummary_l_inst_l_quantity_cmd_ready,
    l_quantity_cmd_firstIdx => PriceSummary_l_inst_l_quantity_cmd_firstIdx,
    l_quantity_cmd_lastIdx => PriceSummary_l_inst_l_quantity_cmd_lastIdx,
    l_quantity_cmd_ctrl => PriceSummary_l_inst_l_quantity_cmd_ctrl,
    l_quantity_cmd_tag => PriceSummary_l_inst_l_quantity_cmd_tag,
    l_quantity_unl_valid => PriceSummary_l_inst_l_quantity_unl_valid,
    l_quantity_unl_ready => PriceSummary_l_inst_l_quantity_unl_ready,
    l_quantity_unl_tag => PriceSummary_l_inst_l_quantity_unl_tag,
    l_extendedprice_valid => PriceSummary_l_inst_l_extendedprice_valid,
    l_extendedprice_ready => PriceSummary_l_inst_l_extendedprice_ready,
    l_extendedprice_dvalid => PriceSummary_l_inst_l_extendedprice_dvalid,
    l_extendedprice_last => PriceSummary_l_inst_l_extendedprice_last,
    l_extendedprice => PriceSummary_l_inst_l_extendedprice,
    l_extendedprice_bus_rreq_valid => PriceSummary_l_inst_l_extendedprice_bus_rreq_valid,
    l_extendedprice_bus_rreq_ready => PriceSummary_l_inst_l_extendedprice_bus_rreq_ready,
    l_extendedprice_bus_rreq_addr => PriceSummary_l_inst_l_extendedprice_bus_rreq_addr,
    l_extendedprice_bus_rreq_len => PriceSummary_l_inst_l_extendedprice_bus_rreq_len,
    l_extendedprice_bus_rdat_valid => PriceSummary_l_inst_l_extendedprice_bus_rdat_valid,
    l_extendedprice_bus_rdat_ready => PriceSummary_l_inst_l_extendedprice_bus_rdat_ready,
    l_extendedprice_bus_rdat_data => PriceSummary_l_inst_l_extendedprice_bus_rdat_data,
    l_extendedprice_bus_rdat_last => PriceSummary_l_inst_l_extendedprice_bus_rdat_last,
    l_extendedprice_cmd_valid => PriceSummary_l_inst_l_extendedprice_cmd_valid,
    l_extendedprice_cmd_ready => PriceSummary_l_inst_l_extendedprice_cmd_ready,
    l_extendedprice_cmd_firstIdx => PriceSummary_l_inst_l_extendedprice_cmd_firstIdx,
    l_extendedprice_cmd_lastIdx => PriceSummary_l_inst_l_extendedprice_cmd_lastIdx,
    l_extendedprice_cmd_ctrl => PriceSummary_l_inst_l_extendedprice_cmd_ctrl,
    l_extendedprice_cmd_tag => PriceSummary_l_inst_l_extendedprice_cmd_tag,
    l_extendedprice_unl_valid => PriceSummary_l_inst_l_extendedprice_unl_valid,
    l_extendedprice_unl_ready => PriceSummary_l_inst_l_extendedprice_unl_ready,
    l_extendedprice_unl_tag => PriceSummary_l_inst_l_extendedprice_unl_tag,
    l_discount_valid => PriceSummary_l_inst_l_discount_valid,
    l_discount_ready => PriceSummary_l_inst_l_discount_ready,
    l_discount_dvalid => PriceSummary_l_inst_l_discount_dvalid,
    l_discount_last => PriceSummary_l_inst_l_discount_last,
    l_discount => PriceSummary_l_inst_l_discount,
    l_discount_bus_rreq_valid => PriceSummary_l_inst_l_discount_bus_rreq_valid,
    l_discount_bus_rreq_ready => PriceSummary_l_inst_l_discount_bus_rreq_ready,
    l_discount_bus_rreq_addr => PriceSummary_l_inst_l_discount_bus_rreq_addr,
    l_discount_bus_rreq_len => PriceSummary_l_inst_l_discount_bus_rreq_len,
    l_discount_bus_rdat_valid => PriceSummary_l_inst_l_discount_bus_rdat_valid,
    l_discount_bus_rdat_ready => PriceSummary_l_inst_l_discount_bus_rdat_ready,
    l_discount_bus_rdat_data => PriceSummary_l_inst_l_discount_bus_rdat_data,
    l_discount_bus_rdat_last => PriceSummary_l_inst_l_discount_bus_rdat_last,
    l_discount_cmd_valid => PriceSummary_l_inst_l_discount_cmd_valid,
    l_discount_cmd_ready => PriceSummary_l_inst_l_discount_cmd_ready,
    l_discount_cmd_firstIdx => PriceSummary_l_inst_l_discount_cmd_firstIdx,
    l_discount_cmd_lastIdx => PriceSummary_l_inst_l_discount_cmd_lastIdx,
    l_discount_cmd_ctrl => PriceSummary_l_inst_l_discount_cmd_ctrl,
    l_discount_cmd_tag => PriceSummary_l_inst_l_discount_cmd_tag,
    l_discount_unl_valid => PriceSummary_l_inst_l_discount_unl_valid,
    l_discount_unl_ready => PriceSummary_l_inst_l_discount_unl_ready,
    l_discount_unl_tag => PriceSummary_l_inst_l_discount_unl_tag,
    l_tax_valid => PriceSummary_l_inst_l_tax_valid,
    l_tax_ready => PriceSummary_l_inst_l_tax_ready,
    l_tax_dvalid => PriceSummary_l_inst_l_tax_dvalid,
    l_tax_last => PriceSummary_l_inst_l_tax_last,
    l_tax => PriceSummary_l_inst_l_tax,
    l_tax_bus_rreq_valid => PriceSummary_l_inst_l_tax_bus_rreq_valid,
    l_tax_bus_rreq_ready => PriceSummary_l_inst_l_tax_bus_rreq_ready,
    l_tax_bus_rreq_addr => PriceSummary_l_inst_l_tax_bus_rreq_addr,
    l_tax_bus_rreq_len => PriceSummary_l_inst_l_tax_bus_rreq_len,
    l_tax_bus_rdat_valid => PriceSummary_l_inst_l_tax_bus_rdat_valid,
    l_tax_bus_rdat_ready => PriceSummary_l_inst_l_tax_bus_rdat_ready,
    l_tax_bus_rdat_data => PriceSummary_l_inst_l_tax_bus_rdat_data,
    l_tax_bus_rdat_last => PriceSummary_l_inst_l_tax_bus_rdat_last,
    l_tax_cmd_valid => PriceSummary_l_inst_l_tax_cmd_valid,
    l_tax_cmd_ready => PriceSummary_l_inst_l_tax_cmd_ready,
    l_tax_cmd_firstIdx => PriceSummary_l_inst_l_tax_cmd_firstIdx,
    l_tax_cmd_lastIdx => PriceSummary_l_inst_l_tax_cmd_lastIdx,
    l_tax_cmd_ctrl => PriceSummary_l_inst_l_tax_cmd_ctrl,
    l_tax_cmd_tag => PriceSummary_l_inst_l_tax_cmd_tag,
    l_tax_unl_valid => PriceSummary_l_inst_l_tax_unl_valid,
    l_tax_unl_ready => PriceSummary_l_inst_l_tax_unl_ready,
    l_tax_unl_tag => PriceSummary_l_inst_l_tax_unl_tag,
    l_returnflag_valid => PriceSummary_l_inst_l_returnflag_valid,
    l_returnflag_ready => PriceSummary_l_inst_l_returnflag_ready,
    l_returnflag_dvalid => PriceSummary_l_inst_l_returnflag_dvalid,
    l_returnflag_last => PriceSummary_l_inst_l_returnflag_last,
    l_returnflag_length => PriceSummary_l_inst_l_returnflag_length,
    l_returnflag_count => PriceSummary_l_inst_l_returnflag_count,
    l_returnflag_chars_valid => PriceSummary_l_inst_l_returnflag_chars_valid,
    l_returnflag_chars_ready => PriceSummary_l_inst_l_returnflag_chars_ready,
    l_returnflag_chars_dvalid => PriceSummary_l_inst_l_returnflag_chars_dvalid,
    l_returnflag_chars_last => PriceSummary_l_inst_l_returnflag_chars_last,
    l_returnflag_chars => PriceSummary_l_inst_l_returnflag_chars,
    l_returnflag_chars_count => PriceSummary_l_inst_l_returnflag_chars_count,
    l_returnflag_bus_rreq_valid => PriceSummary_l_inst_l_returnflag_bus_rreq_valid,
    l_returnflag_bus_rreq_ready => PriceSummary_l_inst_l_returnflag_bus_rreq_ready,
    l_returnflag_bus_rreq_addr => PriceSummary_l_inst_l_returnflag_bus_rreq_addr,
    l_returnflag_bus_rreq_len => PriceSummary_l_inst_l_returnflag_bus_rreq_len,
    l_returnflag_bus_rdat_valid => PriceSummary_l_inst_l_returnflag_bus_rdat_valid,
    l_returnflag_bus_rdat_ready => PriceSummary_l_inst_l_returnflag_bus_rdat_ready,
    l_returnflag_bus_rdat_data => PriceSummary_l_inst_l_returnflag_bus_rdat_data,
    l_returnflag_bus_rdat_last => PriceSummary_l_inst_l_returnflag_bus_rdat_last,
    l_returnflag_cmd_valid => PriceSummary_l_inst_l_returnflag_cmd_valid,
    l_returnflag_cmd_ready => PriceSummary_l_inst_l_returnflag_cmd_ready,
    l_returnflag_cmd_firstIdx => PriceSummary_l_inst_l_returnflag_cmd_firstIdx,
    l_returnflag_cmd_lastIdx => PriceSummary_l_inst_l_returnflag_cmd_lastIdx,
    l_returnflag_cmd_ctrl => PriceSummary_l_inst_l_returnflag_cmd_ctrl,
    l_returnflag_cmd_tag => PriceSummary_l_inst_l_returnflag_cmd_tag,
    l_returnflag_unl_valid => PriceSummary_l_inst_l_returnflag_unl_valid,
    l_returnflag_unl_ready => PriceSummary_l_inst_l_returnflag_unl_ready,
    l_returnflag_unl_tag => PriceSummary_l_inst_l_returnflag_unl_tag,
    l_linestatus_valid => PriceSummary_l_inst_l_linestatus_valid,
    l_linestatus_ready => PriceSummary_l_inst_l_linestatus_ready,
    l_linestatus_dvalid => PriceSummary_l_inst_l_linestatus_dvalid,
    l_linestatus_last => PriceSummary_l_inst_l_linestatus_last,
    l_linestatus_length => PriceSummary_l_inst_l_linestatus_length,
    l_linestatus_count => PriceSummary_l_inst_l_linestatus_count,
    l_linestatus_chars_valid => PriceSummary_l_inst_l_linestatus_chars_valid,
    l_linestatus_chars_ready => PriceSummary_l_inst_l_linestatus_chars_ready,
    l_linestatus_chars_dvalid => PriceSummary_l_inst_l_linestatus_chars_dvalid,
    l_linestatus_chars_last => PriceSummary_l_inst_l_linestatus_chars_last,
    l_linestatus_chars => PriceSummary_l_inst_l_linestatus_chars,
    l_linestatus_chars_count => PriceSummary_l_inst_l_linestatus_chars_count,
    l_linestatus_bus_rreq_valid => PriceSummary_l_inst_l_linestatus_bus_rreq_valid,
    l_linestatus_bus_rreq_ready => PriceSummary_l_inst_l_linestatus_bus_rreq_ready,
    l_linestatus_bus_rreq_addr => PriceSummary_l_inst_l_linestatus_bus_rreq_addr,
    l_linestatus_bus_rreq_len => PriceSummary_l_inst_l_linestatus_bus_rreq_len,
    l_linestatus_bus_rdat_valid => PriceSummary_l_inst_l_linestatus_bus_rdat_valid,
    l_linestatus_bus_rdat_ready => PriceSummary_l_inst_l_linestatus_bus_rdat_ready,
    l_linestatus_bus_rdat_data => PriceSummary_l_inst_l_linestatus_bus_rdat_data,
    l_linestatus_bus_rdat_last => PriceSummary_l_inst_l_linestatus_bus_rdat_last,
    l_linestatus_cmd_valid => PriceSummary_l_inst_l_linestatus_cmd_valid,
    l_linestatus_cmd_ready => PriceSummary_l_inst_l_linestatus_cmd_ready,
    l_linestatus_cmd_firstIdx => PriceSummary_l_inst_l_linestatus_cmd_firstIdx,
    l_linestatus_cmd_lastIdx => PriceSummary_l_inst_l_linestatus_cmd_lastIdx,
    l_linestatus_cmd_ctrl => PriceSummary_l_inst_l_linestatus_cmd_ctrl,
    l_linestatus_cmd_tag => PriceSummary_l_inst_l_linestatus_cmd_tag,
    l_linestatus_unl_valid => PriceSummary_l_inst_l_linestatus_unl_valid,
    l_linestatus_unl_ready => PriceSummary_l_inst_l_linestatus_unl_ready,
    l_linestatus_unl_tag => PriceSummary_l_inst_l_linestatus_unl_tag,
    l_shipdate_valid => PriceSummary_l_inst_l_shipdate_valid,
    l_shipdate_ready => PriceSummary_l_inst_l_shipdate_ready,
    l_shipdate_dvalid => PriceSummary_l_inst_l_shipdate_dvalid,
    l_shipdate_last => PriceSummary_l_inst_l_shipdate_last,
    l_shipdate => PriceSummary_l_inst_l_shipdate,
    l_shipdate_bus_rreq_valid => PriceSummary_l_inst_l_shipdate_bus_rreq_valid,
    l_shipdate_bus_rreq_ready => PriceSummary_l_inst_l_shipdate_bus_rreq_ready,
    l_shipdate_bus_rreq_addr => PriceSummary_l_inst_l_shipdate_bus_rreq_addr,
    l_shipdate_bus_rreq_len => PriceSummary_l_inst_l_shipdate_bus_rreq_len,
    l_shipdate_bus_rdat_valid => PriceSummary_l_inst_l_shipdate_bus_rdat_valid,
    l_shipdate_bus_rdat_ready => PriceSummary_l_inst_l_shipdate_bus_rdat_ready,
    l_shipdate_bus_rdat_data => PriceSummary_l_inst_l_shipdate_bus_rdat_data,
    l_shipdate_bus_rdat_last => PriceSummary_l_inst_l_shipdate_bus_rdat_last,
    l_shipdate_cmd_valid => PriceSummary_l_inst_l_shipdate_cmd_valid,
    l_shipdate_cmd_ready => PriceSummary_l_inst_l_shipdate_cmd_ready,
    l_shipdate_cmd_firstIdx => PriceSummary_l_inst_l_shipdate_cmd_firstIdx,
    l_shipdate_cmd_lastIdx => PriceSummary_l_inst_l_shipdate_cmd_lastIdx,
    l_shipdate_cmd_ctrl => PriceSummary_l_inst_l_shipdate_cmd_ctrl,
    l_shipdate_cmd_tag => PriceSummary_l_inst_l_shipdate_cmd_tag,
    l_shipdate_unl_valid => PriceSummary_l_inst_l_shipdate_unl_valid,
    l_shipdate_unl_ready => PriceSummary_l_inst_l_shipdate_unl_ready,
    l_shipdate_unl_tag => PriceSummary_l_inst_l_shipdate_unl_tag,
    l_returnflag_o_valid => PriceSummaryWriter_l_inst_l_returnflag_o_valid,
    l_returnflag_o_ready => PriceSummaryWriter_l_inst_l_returnflag_o_ready,
    l_returnflag_o_dvalid => PriceSummaryWriter_l_inst_l_returnflag_o_dvalid,
    l_returnflag_o_last => PriceSummaryWriter_l_inst_l_returnflag_o_last,
    l_returnflag_o_length => PriceSummaryWriter_l_inst_l_returnflag_o_length,
    l_returnflag_o_count => PriceSummaryWriter_l_inst_l_returnflag_o_count,
    l_returnflag_o_chars_valid => PriceSummaryWriter_l_inst_l_returnflag_o_chars_valid,
    l_returnflag_o_chars_ready => PriceSummaryWriter_l_inst_l_returnflag_o_chars_ready,
    l_returnflag_o_chars_dvalid => PriceSummaryWriter_l_inst_l_returnflag_o_chars_dvalid,
    l_returnflag_o_chars_last => PriceSummaryWriter_l_inst_l_returnflag_o_chars_last,
    l_returnflag_o_chars => PriceSummaryWriter_l_inst_l_returnflag_o_chars,
    l_returnflag_o_chars_count => PriceSummaryWriter_l_inst_l_returnflag_o_chars_count,
    l_returnflag_o_bus_wreq_valid => PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_valid,
    l_returnflag_o_bus_wreq_ready => PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_ready,
    l_returnflag_o_bus_wreq_addr => PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_addr,
    l_returnflag_o_bus_wreq_len => PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_len,
    l_returnflag_o_bus_wdat_valid => PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_valid,
    l_returnflag_o_bus_wdat_ready => PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_ready,
    l_returnflag_o_bus_wdat_data => PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_data,
    l_returnflag_o_bus_wdat_strobe => PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_strobe,
    l_returnflag_o_bus_wdat_last => PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_last,
    l_returnflag_o_cmd_valid => PriceSummaryWriter_l_inst_l_returnflag_o_cmd_valid,
    l_returnflag_o_cmd_ready => PriceSummaryWriter_l_inst_l_returnflag_o_cmd_ready,
    l_returnflag_o_cmd_firstIdx => PriceSummaryWriter_l_inst_l_returnflag_o_cmd_firstIdx,
    l_returnflag_o_cmd_lastIdx => PriceSummaryWriter_l_inst_l_returnflag_o_cmd_lastIdx,
    l_returnflag_o_cmd_ctrl => PriceSummaryWriter_l_inst_l_returnflag_o_cmd_ctrl,
    l_returnflag_o_cmd_tag => PriceSummaryWriter_l_inst_l_returnflag_o_cmd_tag,
    l_returnflag_o_unl_valid => PriceSummaryWriter_l_inst_l_returnflag_o_unl_valid,
    l_returnflag_o_unl_ready => PriceSummaryWriter_l_inst_l_returnflag_o_unl_ready,
    l_returnflag_o_unl_tag => PriceSummaryWriter_l_inst_l_returnflag_o_unl_tag,
    l_linestatus_o_valid => PriceSummaryWriter_l_inst_l_linestatus_o_valid,
    l_linestatus_o_ready => PriceSummaryWriter_l_inst_l_linestatus_o_ready,
    l_linestatus_o_dvalid => PriceSummaryWriter_l_inst_l_linestatus_o_dvalid,
    l_linestatus_o_last => PriceSummaryWriter_l_inst_l_linestatus_o_last,
    l_linestatus_o_length => PriceSummaryWriter_l_inst_l_linestatus_o_length,
    l_linestatus_o_count => PriceSummaryWriter_l_inst_l_linestatus_o_count,
    l_linestatus_o_chars_valid => PriceSummaryWriter_l_inst_l_linestatus_o_chars_valid,
    l_linestatus_o_chars_ready => PriceSummaryWriter_l_inst_l_linestatus_o_chars_ready,
    l_linestatus_o_chars_dvalid => PriceSummaryWriter_l_inst_l_linestatus_o_chars_dvalid,
    l_linestatus_o_chars_last => PriceSummaryWriter_l_inst_l_linestatus_o_chars_last,
    l_linestatus_o_chars => PriceSummaryWriter_l_inst_l_linestatus_o_chars,
    l_linestatus_o_chars_count => PriceSummaryWriter_l_inst_l_linestatus_o_chars_count,
    l_linestatus_o_bus_wreq_valid => PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_valid,
    l_linestatus_o_bus_wreq_ready => PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_ready,
    l_linestatus_o_bus_wreq_addr => PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_addr,
    l_linestatus_o_bus_wreq_len => PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_len,
    l_linestatus_o_bus_wdat_valid => PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_valid,
    l_linestatus_o_bus_wdat_ready => PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_ready,
    l_linestatus_o_bus_wdat_data => PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_data,
    l_linestatus_o_bus_wdat_strobe => PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_strobe,
    l_linestatus_o_bus_wdat_last => PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_last,
    l_linestatus_o_cmd_valid => PriceSummaryWriter_l_inst_l_linestatus_o_cmd_valid,
    l_linestatus_o_cmd_ready => PriceSummaryWriter_l_inst_l_linestatus_o_cmd_ready,
    l_linestatus_o_cmd_firstIdx => PriceSummaryWriter_l_inst_l_linestatus_o_cmd_firstIdx,
    l_linestatus_o_cmd_lastIdx => PriceSummaryWriter_l_inst_l_linestatus_o_cmd_lastIdx,
    l_linestatus_o_cmd_ctrl => PriceSummaryWriter_l_inst_l_linestatus_o_cmd_ctrl,
    l_linestatus_o_cmd_tag => PriceSummaryWriter_l_inst_l_linestatus_o_cmd_tag,
    l_linestatus_o_unl_valid => PriceSummaryWriter_l_inst_l_linestatus_o_unl_valid,
    l_linestatus_o_unl_ready => PriceSummaryWriter_l_inst_l_linestatus_o_unl_ready,
    l_linestatus_o_unl_tag => PriceSummaryWriter_l_inst_l_linestatus_o_unl_tag,
    l_sum_qty_valid => PriceSummaryWriter_l_inst_l_sum_qty_valid,
    l_sum_qty_ready => PriceSummaryWriter_l_inst_l_sum_qty_ready,
    l_sum_qty_dvalid => PriceSummaryWriter_l_inst_l_sum_qty_dvalid,
    l_sum_qty_last => PriceSummaryWriter_l_inst_l_sum_qty_last,
    l_sum_qty => PriceSummaryWriter_l_inst_l_sum_qty,
    l_sum_qty_bus_wreq_valid => PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_valid,
    l_sum_qty_bus_wreq_ready => PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_ready,
    l_sum_qty_bus_wreq_addr => PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_addr,
    l_sum_qty_bus_wreq_len => PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_len,
    l_sum_qty_bus_wdat_valid => PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_valid,
    l_sum_qty_bus_wdat_ready => PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_ready,
    l_sum_qty_bus_wdat_data => PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_data,
    l_sum_qty_bus_wdat_strobe => PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_strobe,
    l_sum_qty_bus_wdat_last => PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_last,
    l_sum_qty_cmd_valid => PriceSummaryWriter_l_inst_l_sum_qty_cmd_valid,
    l_sum_qty_cmd_ready => PriceSummaryWriter_l_inst_l_sum_qty_cmd_ready,
    l_sum_qty_cmd_firstIdx => PriceSummaryWriter_l_inst_l_sum_qty_cmd_firstIdx,
    l_sum_qty_cmd_lastIdx => PriceSummaryWriter_l_inst_l_sum_qty_cmd_lastIdx,
    l_sum_qty_cmd_ctrl => PriceSummaryWriter_l_inst_l_sum_qty_cmd_ctrl,
    l_sum_qty_cmd_tag => PriceSummaryWriter_l_inst_l_sum_qty_cmd_tag,
    l_sum_qty_unl_valid => PriceSummaryWriter_l_inst_l_sum_qty_unl_valid,
    l_sum_qty_unl_ready => PriceSummaryWriter_l_inst_l_sum_qty_unl_ready,
    l_sum_qty_unl_tag => PriceSummaryWriter_l_inst_l_sum_qty_unl_tag,
    l_sum_base_price_valid => PriceSummaryWriter_l_inst_l_sum_base_price_valid,
    l_sum_base_price_ready => PriceSummaryWriter_l_inst_l_sum_base_price_ready,
    l_sum_base_price_dvalid => PriceSummaryWriter_l_inst_l_sum_base_price_dvalid,
    l_sum_base_price_last => PriceSummaryWriter_l_inst_l_sum_base_price_last,
    l_sum_base_price => PriceSummaryWriter_l_inst_l_sum_base_price,
    l_sum_base_price_bus_wreq_valid => PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_valid,
    l_sum_base_price_bus_wreq_ready => PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_ready,
    l_sum_base_price_bus_wreq_addr => PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_addr,
    l_sum_base_price_bus_wreq_len => PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_len,
    l_sum_base_price_bus_wdat_valid => PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_valid,
    l_sum_base_price_bus_wdat_ready => PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_ready,
    l_sum_base_price_bus_wdat_data => PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_data,
    l_sum_base_price_bus_wdat_strobe => PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_strobe,
    l_sum_base_price_bus_wdat_last => PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_last,
    l_sum_base_price_cmd_valid => PriceSummaryWriter_l_inst_l_sum_base_price_cmd_valid,
    l_sum_base_price_cmd_ready => PriceSummaryWriter_l_inst_l_sum_base_price_cmd_ready,
    l_sum_base_price_cmd_firstIdx => PriceSummaryWriter_l_inst_l_sum_base_price_cmd_firstIdx,
    l_sum_base_price_cmd_lastIdx => PriceSummaryWriter_l_inst_l_sum_base_price_cmd_lastIdx,
    l_sum_base_price_cmd_ctrl => PriceSummaryWriter_l_inst_l_sum_base_price_cmd_ctrl,
    l_sum_base_price_cmd_tag => PriceSummaryWriter_l_inst_l_sum_base_price_cmd_tag,
    l_sum_base_price_unl_valid => PriceSummaryWriter_l_inst_l_sum_base_price_unl_valid,
    l_sum_base_price_unl_ready => PriceSummaryWriter_l_inst_l_sum_base_price_unl_ready,
    l_sum_base_price_unl_tag => PriceSummaryWriter_l_inst_l_sum_base_price_unl_tag,
    l_sum_disc_price_valid => PriceSummaryWriter_l_inst_l_sum_disc_price_valid,
    l_sum_disc_price_ready => PriceSummaryWriter_l_inst_l_sum_disc_price_ready,
    l_sum_disc_price_dvalid => PriceSummaryWriter_l_inst_l_sum_disc_price_dvalid,
    l_sum_disc_price_last => PriceSummaryWriter_l_inst_l_sum_disc_price_last,
    l_sum_disc_price => PriceSummaryWriter_l_inst_l_sum_disc_price,
    l_sum_disc_price_bus_wreq_valid => PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_valid,
    l_sum_disc_price_bus_wreq_ready => PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_ready,
    l_sum_disc_price_bus_wreq_addr => PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_addr,
    l_sum_disc_price_bus_wreq_len => PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_len,
    l_sum_disc_price_bus_wdat_valid => PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_valid,
    l_sum_disc_price_bus_wdat_ready => PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_ready,
    l_sum_disc_price_bus_wdat_data => PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_data,
    l_sum_disc_price_bus_wdat_strobe => PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_strobe,
    l_sum_disc_price_bus_wdat_last => PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_last,
    l_sum_disc_price_cmd_valid => PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_valid,
    l_sum_disc_price_cmd_ready => PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_ready,
    l_sum_disc_price_cmd_firstIdx => PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_firstIdx,
    l_sum_disc_price_cmd_lastIdx => PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_lastIdx,
    l_sum_disc_price_cmd_ctrl => PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_ctrl,
    l_sum_disc_price_cmd_tag => PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_tag,
    l_sum_disc_price_unl_valid => PriceSummaryWriter_l_inst_l_sum_disc_price_unl_valid,
    l_sum_disc_price_unl_ready => PriceSummaryWriter_l_inst_l_sum_disc_price_unl_ready,
    l_sum_disc_price_unl_tag => PriceSummaryWriter_l_inst_l_sum_disc_price_unl_tag,
    l_sum_charge_valid => PriceSummaryWriter_l_inst_l_sum_charge_valid,
    l_sum_charge_ready => PriceSummaryWriter_l_inst_l_sum_charge_ready,
    l_sum_charge_dvalid => PriceSummaryWriter_l_inst_l_sum_charge_dvalid,
    l_sum_charge_last => PriceSummaryWriter_l_inst_l_sum_charge_last,
    l_sum_charge => PriceSummaryWriter_l_inst_l_sum_charge,
    l_sum_charge_bus_wreq_valid => PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_valid,
    l_sum_charge_bus_wreq_ready => PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_ready,
    l_sum_charge_bus_wreq_addr => PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_addr,
    l_sum_charge_bus_wreq_len => PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_len,
    l_sum_charge_bus_wdat_valid => PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_valid,
    l_sum_charge_bus_wdat_ready => PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_ready,
    l_sum_charge_bus_wdat_data => PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_data,
    l_sum_charge_bus_wdat_strobe => PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_strobe,
    l_sum_charge_bus_wdat_last => PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_last,
    l_sum_charge_cmd_valid => PriceSummaryWriter_l_inst_l_sum_charge_cmd_valid,
    l_sum_charge_cmd_ready => PriceSummaryWriter_l_inst_l_sum_charge_cmd_ready,
    l_sum_charge_cmd_firstIdx => PriceSummaryWriter_l_inst_l_sum_charge_cmd_firstIdx,
    l_sum_charge_cmd_lastIdx => PriceSummaryWriter_l_inst_l_sum_charge_cmd_lastIdx,
    l_sum_charge_cmd_ctrl => PriceSummaryWriter_l_inst_l_sum_charge_cmd_ctrl,
    l_sum_charge_cmd_tag => PriceSummaryWriter_l_inst_l_sum_charge_cmd_tag,
    l_sum_charge_unl_valid => PriceSummaryWriter_l_inst_l_sum_charge_unl_valid,
    l_sum_charge_unl_ready => PriceSummaryWriter_l_inst_l_sum_charge_unl_ready,
    l_sum_charge_unl_tag => PriceSummaryWriter_l_inst_l_sum_charge_unl_tag,
    l_avg_qty_valid => PriceSummaryWriter_l_inst_l_avg_qty_valid,
    l_avg_qty_ready => PriceSummaryWriter_l_inst_l_avg_qty_ready,
    l_avg_qty_dvalid => PriceSummaryWriter_l_inst_l_avg_qty_dvalid,
    l_avg_qty_last => PriceSummaryWriter_l_inst_l_avg_qty_last,
    l_avg_qty => PriceSummaryWriter_l_inst_l_avg_qty,
    l_avg_qty_bus_wreq_valid => PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_valid,
    l_avg_qty_bus_wreq_ready => PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_ready,
    l_avg_qty_bus_wreq_addr => PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_addr,
    l_avg_qty_bus_wreq_len => PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_len,
    l_avg_qty_bus_wdat_valid => PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_valid,
    l_avg_qty_bus_wdat_ready => PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_ready,
    l_avg_qty_bus_wdat_data => PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_data,
    l_avg_qty_bus_wdat_strobe => PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_strobe,
    l_avg_qty_bus_wdat_last => PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_last,
    l_avg_qty_cmd_valid => PriceSummaryWriter_l_inst_l_avg_qty_cmd_valid,
    l_avg_qty_cmd_ready => PriceSummaryWriter_l_inst_l_avg_qty_cmd_ready,
    l_avg_qty_cmd_firstIdx => PriceSummaryWriter_l_inst_l_avg_qty_cmd_firstIdx,
    l_avg_qty_cmd_lastIdx => PriceSummaryWriter_l_inst_l_avg_qty_cmd_lastIdx,
    l_avg_qty_cmd_ctrl => PriceSummaryWriter_l_inst_l_avg_qty_cmd_ctrl,
    l_avg_qty_cmd_tag => PriceSummaryWriter_l_inst_l_avg_qty_cmd_tag,
    l_avg_qty_unl_valid => PriceSummaryWriter_l_inst_l_avg_qty_unl_valid,
    l_avg_qty_unl_ready => PriceSummaryWriter_l_inst_l_avg_qty_unl_ready,
    l_avg_qty_unl_tag => PriceSummaryWriter_l_inst_l_avg_qty_unl_tag,
    l_avg_price_valid => PriceSummaryWriter_l_inst_l_avg_price_valid,
    l_avg_price_ready => PriceSummaryWriter_l_inst_l_avg_price_ready,
    l_avg_price_dvalid => PriceSummaryWriter_l_inst_l_avg_price_dvalid,
    l_avg_price_last => PriceSummaryWriter_l_inst_l_avg_price_last,
    l_avg_price => PriceSummaryWriter_l_inst_l_avg_price,
    l_avg_price_bus_wreq_valid => PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_valid,
    l_avg_price_bus_wreq_ready => PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_ready,
    l_avg_price_bus_wreq_addr => PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_addr,
    l_avg_price_bus_wreq_len => PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_len,
    l_avg_price_bus_wdat_valid => PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_valid,
    l_avg_price_bus_wdat_ready => PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_ready,
    l_avg_price_bus_wdat_data => PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_data,
    l_avg_price_bus_wdat_strobe => PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_strobe,
    l_avg_price_bus_wdat_last => PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_last,
    l_avg_price_cmd_valid => PriceSummaryWriter_l_inst_l_avg_price_cmd_valid,
    l_avg_price_cmd_ready => PriceSummaryWriter_l_inst_l_avg_price_cmd_ready,
    l_avg_price_cmd_firstIdx => PriceSummaryWriter_l_inst_l_avg_price_cmd_firstIdx,
    l_avg_price_cmd_lastIdx => PriceSummaryWriter_l_inst_l_avg_price_cmd_lastIdx,
    l_avg_price_cmd_ctrl => PriceSummaryWriter_l_inst_l_avg_price_cmd_ctrl,
    l_avg_price_cmd_tag => PriceSummaryWriter_l_inst_l_avg_price_cmd_tag,
    l_avg_price_unl_valid => PriceSummaryWriter_l_inst_l_avg_price_unl_valid,
    l_avg_price_unl_ready => PriceSummaryWriter_l_inst_l_avg_price_unl_ready,
    l_avg_price_unl_tag => PriceSummaryWriter_l_inst_l_avg_price_unl_tag,
    l_avg_disc_valid => PriceSummaryWriter_l_inst_l_avg_disc_valid,
    l_avg_disc_ready => PriceSummaryWriter_l_inst_l_avg_disc_ready,
    l_avg_disc_dvalid => PriceSummaryWriter_l_inst_l_avg_disc_dvalid,
    l_avg_disc_last => PriceSummaryWriter_l_inst_l_avg_disc_last,
    l_avg_disc => PriceSummaryWriter_l_inst_l_avg_disc,
    l_avg_disc_bus_wreq_valid => PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_valid,
    l_avg_disc_bus_wreq_ready => PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_ready,
    l_avg_disc_bus_wreq_addr => PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_addr,
    l_avg_disc_bus_wreq_len => PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_len,
    l_avg_disc_bus_wdat_valid => PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_valid,
    l_avg_disc_bus_wdat_ready => PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_ready,
    l_avg_disc_bus_wdat_data => PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_data,
    l_avg_disc_bus_wdat_strobe => PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_strobe,
    l_avg_disc_bus_wdat_last => PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_last,
    l_avg_disc_cmd_valid => PriceSummaryWriter_l_inst_l_avg_disc_cmd_valid,
    l_avg_disc_cmd_ready => PriceSummaryWriter_l_inst_l_avg_disc_cmd_ready,
    l_avg_disc_cmd_firstIdx => PriceSummaryWriter_l_inst_l_avg_disc_cmd_firstIdx,
    l_avg_disc_cmd_lastIdx => PriceSummaryWriter_l_inst_l_avg_disc_cmd_lastIdx,
    l_avg_disc_cmd_ctrl => PriceSummaryWriter_l_inst_l_avg_disc_cmd_ctrl,
    l_avg_disc_cmd_tag => PriceSummaryWriter_l_inst_l_avg_disc_cmd_tag,
    l_avg_disc_unl_valid => PriceSummaryWriter_l_inst_l_avg_disc_unl_valid,
    l_avg_disc_unl_ready => PriceSummaryWriter_l_inst_l_avg_disc_unl_ready,
    l_avg_disc_unl_tag => PriceSummaryWriter_l_inst_l_avg_disc_unl_tag,
    l_count_order_valid => PriceSummaryWriter_l_inst_l_count_order_valid,
    l_count_order_ready => PriceSummaryWriter_l_inst_l_count_order_ready,
    l_count_order_dvalid => PriceSummaryWriter_l_inst_l_count_order_dvalid,
    l_count_order_last => PriceSummaryWriter_l_inst_l_count_order_last,
    l_count_order => PriceSummaryWriter_l_inst_l_count_order,
    l_count_order_bus_wreq_valid => PriceSummaryWriter_l_inst_l_count_order_bus_wreq_valid,
    l_count_order_bus_wreq_ready => PriceSummaryWriter_l_inst_l_count_order_bus_wreq_ready,
    l_count_order_bus_wreq_addr => PriceSummaryWriter_l_inst_l_count_order_bus_wreq_addr,
    l_count_order_bus_wreq_len => PriceSummaryWriter_l_inst_l_count_order_bus_wreq_len,
    l_count_order_bus_wdat_valid => PriceSummaryWriter_l_inst_l_count_order_bus_wdat_valid,
    l_count_order_bus_wdat_ready => PriceSummaryWriter_l_inst_l_count_order_bus_wdat_ready,
    l_count_order_bus_wdat_data => PriceSummaryWriter_l_inst_l_count_order_bus_wdat_data,
    l_count_order_bus_wdat_strobe => PriceSummaryWriter_l_inst_l_count_order_bus_wdat_strobe,
    l_count_order_bus_wdat_last => PriceSummaryWriter_l_inst_l_count_order_bus_wdat_last,
    l_count_order_cmd_valid => PriceSummaryWriter_l_inst_l_count_order_cmd_valid,
    l_count_order_cmd_ready => PriceSummaryWriter_l_inst_l_count_order_cmd_ready,
    l_count_order_cmd_firstIdx => PriceSummaryWriter_l_inst_l_count_order_cmd_firstIdx,
    l_count_order_cmd_lastIdx => PriceSummaryWriter_l_inst_l_count_order_cmd_lastIdx,
    l_count_order_cmd_ctrl => PriceSummaryWriter_l_inst_l_count_order_cmd_ctrl,
    l_count_order_cmd_tag => PriceSummaryWriter_l_inst_l_count_order_cmd_tag,
    l_count_order_unl_valid => PriceSummaryWriter_l_inst_l_count_order_unl_valid,
    l_count_order_unl_ready => PriceSummaryWriter_l_inst_l_count_order_unl_ready,
    l_count_order_unl_tag => PriceSummaryWriter_l_inst_l_count_order_unl_tag
  );

  WRAW64DW512LW8BS1BM16_inst : BusWriteArbiterVec
  GENERIC MAP(
    BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    BUS_DATA_WIDTH => BUS_DATA_WIDTH,
    BUS_LEN_WIDTH => BUS_LEN_WIDTH,
    NUM_SLAVE_PORTS => 10,
    ARB_METHOD => "RR-STICKY",
    MAX_OUTSTANDING => 4,
    RAM_CONFIG => "",
    SLV_REQ_SLICES => true,
    MST_REQ_SLICE => true,
    MST_DAT_SLICE => true,
    SLV_DAT_SLICES => true
  )
  PORT MAP(
    bcd_clk => bcd_clk,
    bcd_reset => bcd_reset,
    mst_wreq_valid => WRAW64DW512LW8BS1BM16_inst_mst_wreq_valid,
    mst_wreq_ready => WRAW64DW512LW8BS1BM16_inst_mst_wreq_ready,
    mst_wreq_addr => WRAW64DW512LW8BS1BM16_inst_mst_wreq_addr,
    mst_wreq_len => WRAW64DW512LW8BS1BM16_inst_mst_wreq_len,
    mst_wdat_valid => WRAW64DW512LW8BS1BM16_inst_mst_wdat_valid,
    mst_wdat_ready => WRAW64DW512LW8BS1BM16_inst_mst_wdat_ready,
    mst_wdat_data => WRAW64DW512LW8BS1BM16_inst_mst_wdat_data,
    mst_wdat_strobe => WRAW64DW512LW8BS1BM16_inst_mst_wdat_strobe,
    mst_wdat_last => WRAW64DW512LW8BS1BM16_inst_mst_wdat_last,
    bsv_wreq_valid => WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid,
    bsv_wreq_ready => WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready,
    bsv_wreq_len => WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len,
    bsv_wreq_addr => WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr,
    bsv_wdat_valid => WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid,
    bsv_wdat_strobe => WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe,
    bsv_wdat_ready => WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready,
    bsv_wdat_last => WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last,
    bsv_wdat_data => WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data
  );

  wr_mst_wreq_valid <= WRAW64DW512LW8BS1BM16_inst_mst_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_mst_wreq_ready <= wr_mst_wreq_ready;
  wr_mst_wreq_addr <= WRAW64DW512LW8BS1BM16_inst_mst_wreq_addr;
  wr_mst_wreq_len <= WRAW64DW512LW8BS1BM16_inst_mst_wreq_len;
  wr_mst_wdat_valid <= WRAW64DW512LW8BS1BM16_inst_mst_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_mst_wdat_ready <= wr_mst_wdat_ready;
  wr_mst_wdat_data <= WRAW64DW512LW8BS1BM16_inst_mst_wdat_data;
  wr_mst_wdat_strobe <= WRAW64DW512LW8BS1BM16_inst_mst_wdat_strobe;
  wr_mst_wdat_last <= WRAW64DW512LW8BS1BM16_inst_mst_wdat_last;

  PriceSummaryWriter_Nucleus_inst_l_returnflag_o_unl_valid <= PriceSummaryWriter_l_inst_l_returnflag_o_unl_valid;
  PriceSummaryWriter_l_inst_l_returnflag_o_unl_ready <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_unl_ready;
  PriceSummaryWriter_Nucleus_inst_l_returnflag_o_unl_tag <= PriceSummaryWriter_l_inst_l_returnflag_o_unl_tag;

  PriceSummaryWriter_Nucleus_inst_l_linestatus_o_unl_valid <= PriceSummaryWriter_l_inst_l_linestatus_o_unl_valid;
  PriceSummaryWriter_l_inst_l_linestatus_o_unl_ready <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_unl_ready;
  PriceSummaryWriter_Nucleus_inst_l_linestatus_o_unl_tag <= PriceSummaryWriter_l_inst_l_linestatus_o_unl_tag;

  PriceSummaryWriter_Nucleus_inst_l_sum_qty_unl_valid <= PriceSummaryWriter_l_inst_l_sum_qty_unl_valid;
  PriceSummaryWriter_l_inst_l_sum_qty_unl_ready <= PriceSummaryWriter_Nucleus_inst_l_sum_qty_unl_ready;
  PriceSummaryWriter_Nucleus_inst_l_sum_qty_unl_tag <= PriceSummaryWriter_l_inst_l_sum_qty_unl_tag;

  PriceSummaryWriter_Nucleus_inst_l_sum_base_price_unl_valid <= PriceSummaryWriter_l_inst_l_sum_base_price_unl_valid;
  PriceSummaryWriter_l_inst_l_sum_base_price_unl_ready <= PriceSummaryWriter_Nucleus_inst_l_sum_base_price_unl_ready;
  PriceSummaryWriter_Nucleus_inst_l_sum_base_price_unl_tag <= PriceSummaryWriter_l_inst_l_sum_base_price_unl_tag;

  PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_unl_valid <= PriceSummaryWriter_l_inst_l_sum_disc_price_unl_valid;
  PriceSummaryWriter_l_inst_l_sum_disc_price_unl_ready <= PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_unl_ready;
  PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_unl_tag <= PriceSummaryWriter_l_inst_l_sum_disc_price_unl_tag;

  PriceSummaryWriter_Nucleus_inst_l_sum_charge_unl_valid <= PriceSummaryWriter_l_inst_l_sum_charge_unl_valid;
  PriceSummaryWriter_l_inst_l_sum_charge_unl_ready <= PriceSummaryWriter_Nucleus_inst_l_sum_charge_unl_ready;
  PriceSummaryWriter_Nucleus_inst_l_sum_charge_unl_tag <= PriceSummaryWriter_l_inst_l_sum_charge_unl_tag;

  PriceSummaryWriter_Nucleus_inst_l_avg_qty_unl_valid <= PriceSummaryWriter_l_inst_l_avg_qty_unl_valid;
  PriceSummaryWriter_l_inst_l_avg_qty_unl_ready <= PriceSummaryWriter_Nucleus_inst_l_avg_qty_unl_ready;
  PriceSummaryWriter_Nucleus_inst_l_avg_qty_unl_tag <= PriceSummaryWriter_l_inst_l_avg_qty_unl_tag;

  PriceSummaryWriter_Nucleus_inst_l_avg_price_unl_valid <= PriceSummaryWriter_l_inst_l_avg_price_unl_valid;
  PriceSummaryWriter_l_inst_l_avg_price_unl_ready <= PriceSummaryWriter_Nucleus_inst_l_avg_price_unl_ready;
  PriceSummaryWriter_Nucleus_inst_l_avg_price_unl_tag <= PriceSummaryWriter_l_inst_l_avg_price_unl_tag;

  PriceSummaryWriter_Nucleus_inst_l_avg_disc_unl_valid <= PriceSummaryWriter_l_inst_l_avg_disc_unl_valid;
  PriceSummaryWriter_l_inst_l_avg_disc_unl_ready <= PriceSummaryWriter_Nucleus_inst_l_avg_disc_unl_ready;
  PriceSummaryWriter_Nucleus_inst_l_avg_disc_unl_tag <= PriceSummaryWriter_l_inst_l_avg_disc_unl_tag;

  PriceSummaryWriter_Nucleus_inst_l_count_order_unl_valid <= PriceSummaryWriter_l_inst_l_count_order_unl_valid;
  PriceSummaryWriter_l_inst_l_count_order_unl_ready <= PriceSummaryWriter_Nucleus_inst_l_count_order_unl_ready;
  PriceSummaryWriter_Nucleus_inst_l_count_order_unl_tag <= PriceSummaryWriter_l_inst_l_count_order_unl_tag;

  PriceSummaryWriter_l_inst_l_returnflag_o_valid <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_valid;
  PriceSummaryWriter_Nucleus_inst_l_returnflag_o_ready <= PriceSummaryWriter_l_inst_l_returnflag_o_ready;
  PriceSummaryWriter_l_inst_l_returnflag_o_dvalid <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_dvalid;
  PriceSummaryWriter_l_inst_l_returnflag_o_last <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_last;
  PriceSummaryWriter_l_inst_l_returnflag_o_length <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_length;
  PriceSummaryWriter_l_inst_l_returnflag_o_count <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_count;
  PriceSummaryWriter_l_inst_l_returnflag_o_chars_valid <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_valid;
  PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_ready <= PriceSummaryWriter_l_inst_l_returnflag_o_chars_ready;
  PriceSummaryWriter_l_inst_l_returnflag_o_chars_dvalid <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_dvalid;
  PriceSummaryWriter_l_inst_l_returnflag_o_chars_last <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_last;
  PriceSummaryWriter_l_inst_l_returnflag_o_chars <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars;
  PriceSummaryWriter_l_inst_l_returnflag_o_chars_count <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_count;

  PriceSummaryWriter_l_inst_l_returnflag_o_cmd_valid <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_valid;
  PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_ready <= PriceSummaryWriter_l_inst_l_returnflag_o_cmd_ready;
  PriceSummaryWriter_l_inst_l_returnflag_o_cmd_firstIdx <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_firstIdx;
  PriceSummaryWriter_l_inst_l_returnflag_o_cmd_lastIdx <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_lastIdx;
  PriceSummaryWriter_l_inst_l_returnflag_o_cmd_ctrl <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_ctrl;
  PriceSummaryWriter_l_inst_l_returnflag_o_cmd_tag <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_tag;

  PriceSummaryWriter_l_inst_l_linestatus_o_valid <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_valid;
  PriceSummaryWriter_Nucleus_inst_l_linestatus_o_ready <= PriceSummaryWriter_l_inst_l_linestatus_o_ready;
  PriceSummaryWriter_l_inst_l_linestatus_o_dvalid <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_dvalid;
  PriceSummaryWriter_l_inst_l_linestatus_o_last <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_last;
  PriceSummaryWriter_l_inst_l_linestatus_o_length <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_length;
  PriceSummaryWriter_l_inst_l_linestatus_o_count <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_count;
  PriceSummaryWriter_l_inst_l_linestatus_o_chars_valid <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_valid;
  PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_ready <= PriceSummaryWriter_l_inst_l_linestatus_o_chars_ready;
  PriceSummaryWriter_l_inst_l_linestatus_o_chars_dvalid <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_dvalid;
  PriceSummaryWriter_l_inst_l_linestatus_o_chars_last <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_last;
  PriceSummaryWriter_l_inst_l_linestatus_o_chars <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars;
  PriceSummaryWriter_l_inst_l_linestatus_o_chars_count <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_count;

  PriceSummaryWriter_l_inst_l_linestatus_o_cmd_valid <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_valid;
  PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_ready <= PriceSummaryWriter_l_inst_l_linestatus_o_cmd_ready;
  PriceSummaryWriter_l_inst_l_linestatus_o_cmd_firstIdx <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_firstIdx;
  PriceSummaryWriter_l_inst_l_linestatus_o_cmd_lastIdx <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_lastIdx;
  PriceSummaryWriter_l_inst_l_linestatus_o_cmd_ctrl <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_ctrl;
  PriceSummaryWriter_l_inst_l_linestatus_o_cmd_tag <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_tag;

  PriceSummaryWriter_l_inst_l_sum_qty_valid <= PriceSummaryWriter_Nucleus_inst_l_sum_qty_valid;
  PriceSummaryWriter_Nucleus_inst_l_sum_qty_ready <= PriceSummaryWriter_l_inst_l_sum_qty_ready;
  PriceSummaryWriter_l_inst_l_sum_qty_dvalid <= PriceSummaryWriter_Nucleus_inst_l_sum_qty_dvalid;
  PriceSummaryWriter_l_inst_l_sum_qty_last <= PriceSummaryWriter_Nucleus_inst_l_sum_qty_last;
  PriceSummaryWriter_l_inst_l_sum_qty <= PriceSummaryWriter_Nucleus_inst_l_sum_qty;

  PriceSummaryWriter_l_inst_l_sum_qty_cmd_valid <= PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_valid;
  PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_ready <= PriceSummaryWriter_l_inst_l_sum_qty_cmd_ready;
  PriceSummaryWriter_l_inst_l_sum_qty_cmd_firstIdx <= PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_firstIdx;
  PriceSummaryWriter_l_inst_l_sum_qty_cmd_lastIdx <= PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_lastIdx;
  PriceSummaryWriter_l_inst_l_sum_qty_cmd_ctrl <= PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_ctrl;
  PriceSummaryWriter_l_inst_l_sum_qty_cmd_tag <= PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_tag;

  PriceSummaryWriter_l_inst_l_sum_base_price_valid <= PriceSummaryWriter_Nucleus_inst_l_sum_base_price_valid;
  PriceSummaryWriter_Nucleus_inst_l_sum_base_price_ready <= PriceSummaryWriter_l_inst_l_sum_base_price_ready;
  PriceSummaryWriter_l_inst_l_sum_base_price_dvalid <= PriceSummaryWriter_Nucleus_inst_l_sum_base_price_dvalid;
  PriceSummaryWriter_l_inst_l_sum_base_price_last <= PriceSummaryWriter_Nucleus_inst_l_sum_base_price_last;
  PriceSummaryWriter_l_inst_l_sum_base_price <= PriceSummaryWriter_Nucleus_inst_l_sum_base_price;

  PriceSummaryWriter_l_inst_l_sum_base_price_cmd_valid <= PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_valid;
  PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_ready <= PriceSummaryWriter_l_inst_l_sum_base_price_cmd_ready;
  PriceSummaryWriter_l_inst_l_sum_base_price_cmd_firstIdx <= PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_firstIdx;
  PriceSummaryWriter_l_inst_l_sum_base_price_cmd_lastIdx <= PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_lastIdx;
  PriceSummaryWriter_l_inst_l_sum_base_price_cmd_ctrl <= PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_ctrl;
  PriceSummaryWriter_l_inst_l_sum_base_price_cmd_tag <= PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_tag;

  PriceSummaryWriter_l_inst_l_sum_disc_price_valid <= PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_valid;
  PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_ready <= PriceSummaryWriter_l_inst_l_sum_disc_price_ready;
  PriceSummaryWriter_l_inst_l_sum_disc_price_dvalid <= PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_dvalid;
  PriceSummaryWriter_l_inst_l_sum_disc_price_last <= PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_last;
  PriceSummaryWriter_l_inst_l_sum_disc_price <= PriceSummaryWriter_Nucleus_inst_l_sum_disc_price;

  PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_valid <= PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_valid;
  PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_ready <= PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_ready;
  PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_firstIdx <= PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_firstIdx;
  PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_lastIdx <= PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_lastIdx;
  PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_ctrl <= PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_ctrl;
  PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_tag <= PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_tag;

  PriceSummaryWriter_l_inst_l_sum_charge_valid <= PriceSummaryWriter_Nucleus_inst_l_sum_charge_valid;
  PriceSummaryWriter_Nucleus_inst_l_sum_charge_ready <= PriceSummaryWriter_l_inst_l_sum_charge_ready;
  PriceSummaryWriter_l_inst_l_sum_charge_dvalid <= PriceSummaryWriter_Nucleus_inst_l_sum_charge_dvalid;
  PriceSummaryWriter_l_inst_l_sum_charge_last <= PriceSummaryWriter_Nucleus_inst_l_sum_charge_last;
  PriceSummaryWriter_l_inst_l_sum_charge <= PriceSummaryWriter_Nucleus_inst_l_sum_charge;

  PriceSummaryWriter_l_inst_l_sum_charge_cmd_valid <= PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_valid;
  PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_ready <= PriceSummaryWriter_l_inst_l_sum_charge_cmd_ready;
  PriceSummaryWriter_l_inst_l_sum_charge_cmd_firstIdx <= PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_firstIdx;
  PriceSummaryWriter_l_inst_l_sum_charge_cmd_lastIdx <= PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_lastIdx;
  PriceSummaryWriter_l_inst_l_sum_charge_cmd_ctrl <= PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_ctrl;
  PriceSummaryWriter_l_inst_l_sum_charge_cmd_tag <= PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_tag;

  PriceSummaryWriter_l_inst_l_avg_qty_valid <= PriceSummaryWriter_Nucleus_inst_l_avg_qty_valid;
  PriceSummaryWriter_Nucleus_inst_l_avg_qty_ready <= PriceSummaryWriter_l_inst_l_avg_qty_ready;
  PriceSummaryWriter_l_inst_l_avg_qty_dvalid <= PriceSummaryWriter_Nucleus_inst_l_avg_qty_dvalid;
  PriceSummaryWriter_l_inst_l_avg_qty_last <= PriceSummaryWriter_Nucleus_inst_l_avg_qty_last;
  PriceSummaryWriter_l_inst_l_avg_qty <= PriceSummaryWriter_Nucleus_inst_l_avg_qty;

  PriceSummaryWriter_l_inst_l_avg_qty_cmd_valid <= PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_valid;
  PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_ready <= PriceSummaryWriter_l_inst_l_avg_qty_cmd_ready;
  PriceSummaryWriter_l_inst_l_avg_qty_cmd_firstIdx <= PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_firstIdx;
  PriceSummaryWriter_l_inst_l_avg_qty_cmd_lastIdx <= PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_lastIdx;
  PriceSummaryWriter_l_inst_l_avg_qty_cmd_ctrl <= PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_ctrl;
  PriceSummaryWriter_l_inst_l_avg_qty_cmd_tag <= PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_tag;

  PriceSummaryWriter_l_inst_l_avg_price_valid <= PriceSummaryWriter_Nucleus_inst_l_avg_price_valid;
  PriceSummaryWriter_Nucleus_inst_l_avg_price_ready <= PriceSummaryWriter_l_inst_l_avg_price_ready;
  PriceSummaryWriter_l_inst_l_avg_price_dvalid <= PriceSummaryWriter_Nucleus_inst_l_avg_price_dvalid;
  PriceSummaryWriter_l_inst_l_avg_price_last <= PriceSummaryWriter_Nucleus_inst_l_avg_price_last;
  PriceSummaryWriter_l_inst_l_avg_price <= PriceSummaryWriter_Nucleus_inst_l_avg_price;

  PriceSummaryWriter_l_inst_l_avg_price_cmd_valid <= PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_valid;
  PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_ready <= PriceSummaryWriter_l_inst_l_avg_price_cmd_ready;
  PriceSummaryWriter_l_inst_l_avg_price_cmd_firstIdx <= PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_firstIdx;
  PriceSummaryWriter_l_inst_l_avg_price_cmd_lastIdx <= PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_lastIdx;
  PriceSummaryWriter_l_inst_l_avg_price_cmd_ctrl <= PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_ctrl;
  PriceSummaryWriter_l_inst_l_avg_price_cmd_tag <= PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_tag;

  PriceSummaryWriter_l_inst_l_avg_disc_valid <= PriceSummaryWriter_Nucleus_inst_l_avg_disc_valid;
  PriceSummaryWriter_Nucleus_inst_l_avg_disc_ready <= PriceSummaryWriter_l_inst_l_avg_disc_ready;
  PriceSummaryWriter_l_inst_l_avg_disc_dvalid <= PriceSummaryWriter_Nucleus_inst_l_avg_disc_dvalid;
  PriceSummaryWriter_l_inst_l_avg_disc_last <= PriceSummaryWriter_Nucleus_inst_l_avg_disc_last;
  PriceSummaryWriter_l_inst_l_avg_disc <= PriceSummaryWriter_Nucleus_inst_l_avg_disc;

  PriceSummaryWriter_l_inst_l_avg_disc_cmd_valid <= PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_valid;
  PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_ready <= PriceSummaryWriter_l_inst_l_avg_disc_cmd_ready;
  PriceSummaryWriter_l_inst_l_avg_disc_cmd_firstIdx <= PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_firstIdx;
  PriceSummaryWriter_l_inst_l_avg_disc_cmd_lastIdx <= PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_lastIdx;
  PriceSummaryWriter_l_inst_l_avg_disc_cmd_ctrl <= PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_ctrl;
  PriceSummaryWriter_l_inst_l_avg_disc_cmd_tag <= PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_tag;

  PriceSummaryWriter_l_inst_l_count_order_valid <= PriceSummaryWriter_Nucleus_inst_l_count_order_valid;
  PriceSummaryWriter_Nucleus_inst_l_count_order_ready <= PriceSummaryWriter_l_inst_l_count_order_ready;
  PriceSummaryWriter_l_inst_l_count_order_dvalid <= PriceSummaryWriter_Nucleus_inst_l_count_order_dvalid;
  PriceSummaryWriter_l_inst_l_count_order_last <= PriceSummaryWriter_Nucleus_inst_l_count_order_last;
  PriceSummaryWriter_l_inst_l_count_order <= PriceSummaryWriter_Nucleus_inst_l_count_order;

  PriceSummaryWriter_l_inst_l_count_order_cmd_valid <= PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_valid;
  PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_ready <= PriceSummaryWriter_l_inst_l_count_order_cmd_ready;
  PriceSummaryWriter_l_inst_l_count_order_cmd_firstIdx <= PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_firstIdx;
  PriceSummaryWriter_l_inst_l_count_order_cmd_lastIdx <= PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_lastIdx;
  PriceSummaryWriter_l_inst_l_count_order_cmd_ctrl <= PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_ctrl;
  PriceSummaryWriter_l_inst_l_count_order_cmd_tag <= PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_tag;

  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid(0) <= PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid(1) <= PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid(2) <= PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid(3) <= PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid(4) <= PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid(5) <= PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid(6) <= PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid(7) <= PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid(8) <= PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid(9) <= PriceSummaryWriter_l_inst_l_count_order_bus_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len(BUS_LEN_WIDTH - 1 DOWNTO 0) <= PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_len;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len(BUS_LEN_WIDTH + BUS_LEN_WIDTH - 1 DOWNTO BUS_LEN_WIDTH) <= PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_len;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len(BUS_LEN_WIDTH * 2 + BUS_LEN_WIDTH - 1 DOWNTO BUS_LEN_WIDTH * 2) <= PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_len;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len(BUS_LEN_WIDTH * 3 + BUS_LEN_WIDTH - 1 DOWNTO BUS_LEN_WIDTH * 3) <= PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_len;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len(BUS_LEN_WIDTH * 4 + BUS_LEN_WIDTH - 1 DOWNTO BUS_LEN_WIDTH * 4) <= PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_len;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len(BUS_LEN_WIDTH * 5 + BUS_LEN_WIDTH - 1 DOWNTO BUS_LEN_WIDTH * 5) <= PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_len;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len(BUS_LEN_WIDTH * 6 + BUS_LEN_WIDTH - 1 DOWNTO BUS_LEN_WIDTH * 6) <= PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_len;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len(BUS_LEN_WIDTH * 7 + BUS_LEN_WIDTH - 1 DOWNTO BUS_LEN_WIDTH * 7) <= PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_len;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len(BUS_LEN_WIDTH * 8 + BUS_LEN_WIDTH - 1 DOWNTO BUS_LEN_WIDTH * 8) <= PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_len;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len(BUS_LEN_WIDTH * 9 + BUS_LEN_WIDTH - 1 DOWNTO BUS_LEN_WIDTH * 9) <= PriceSummaryWriter_l_inst_l_count_order_bus_wreq_len;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr(BUS_ADDR_WIDTH - 1 DOWNTO 0) <= PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_addr;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr(BUS_ADDR_WIDTH + BUS_ADDR_WIDTH - 1 DOWNTO BUS_ADDR_WIDTH) <= PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_addr;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr(BUS_ADDR_WIDTH * 2 + BUS_ADDR_WIDTH - 1 DOWNTO BUS_ADDR_WIDTH * 2) <= PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_addr;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr(BUS_ADDR_WIDTH * 3 + BUS_ADDR_WIDTH - 1 DOWNTO BUS_ADDR_WIDTH * 3) <= PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_addr;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr(BUS_ADDR_WIDTH * 4 + BUS_ADDR_WIDTH - 1 DOWNTO BUS_ADDR_WIDTH * 4) <= PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_addr;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr(BUS_ADDR_WIDTH * 5 + BUS_ADDR_WIDTH - 1 DOWNTO BUS_ADDR_WIDTH * 5) <= PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_addr;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr(BUS_ADDR_WIDTH * 6 + BUS_ADDR_WIDTH - 1 DOWNTO BUS_ADDR_WIDTH * 6) <= PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_addr;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr(BUS_ADDR_WIDTH * 7 + BUS_ADDR_WIDTH - 1 DOWNTO BUS_ADDR_WIDTH * 7) <= PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_addr;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr(BUS_ADDR_WIDTH * 8 + BUS_ADDR_WIDTH - 1 DOWNTO BUS_ADDR_WIDTH * 8) <= PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_addr;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr(BUS_ADDR_WIDTH * 9 + BUS_ADDR_WIDTH - 1 DOWNTO BUS_ADDR_WIDTH * 9) <= PriceSummaryWriter_l_inst_l_count_order_bus_wreq_addr;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid(0) <= PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid(1) <= PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid(2) <= PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid(3) <= PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid(4) <= PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid(5) <= PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid(6) <= PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid(7) <= PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid(8) <= PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid(9) <= PriceSummaryWriter_l_inst_l_count_order_bus_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe(BUS_DATA_WIDTH/8 - 1 DOWNTO 0) <= PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_strobe;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe(BUS_DATA_WIDTH/8 + BUS_DATA_WIDTH/8 - 1 DOWNTO BUS_DATA_WIDTH/8) <= PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_strobe;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe(BUS_DATA_WIDTH/8 * 2 + BUS_DATA_WIDTH/8 - 1 DOWNTO BUS_DATA_WIDTH/8 * 2) <= PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_strobe;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe(BUS_DATA_WIDTH/8 * 3 + BUS_DATA_WIDTH/8 - 1 DOWNTO BUS_DATA_WIDTH/8 * 3) <= PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_strobe;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe(BUS_DATA_WIDTH/8 * 4 + BUS_DATA_WIDTH/8 - 1 DOWNTO BUS_DATA_WIDTH/8 * 4) <= PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_strobe;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe(BUS_DATA_WIDTH/8 * 5 + BUS_DATA_WIDTH/8 - 1 DOWNTO BUS_DATA_WIDTH/8 * 5) <= PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_strobe;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe(BUS_DATA_WIDTH/8 * 6 + BUS_DATA_WIDTH/8 - 1 DOWNTO BUS_DATA_WIDTH/8 * 6) <= PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_strobe;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe(BUS_DATA_WIDTH/8 * 7 + BUS_DATA_WIDTH/8 - 1 DOWNTO BUS_DATA_WIDTH/8 * 7) <= PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_strobe;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe(BUS_DATA_WIDTH/8 * 8 + BUS_DATA_WIDTH/8 - 1 DOWNTO BUS_DATA_WIDTH/8 * 8) <= PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_strobe;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe(BUS_DATA_WIDTH/8 * 9 + BUS_DATA_WIDTH/8 - 1 DOWNTO BUS_DATA_WIDTH/8 * 9) <= PriceSummaryWriter_l_inst_l_count_order_bus_wdat_strobe;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last(0) <= PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_last;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last(1) <= PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_last;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last(2) <= PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_last;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last(3) <= PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_last;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last(4) <= PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_last;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last(5) <= PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_last;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last(6) <= PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_last;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last(7) <= PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_last;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last(8) <= PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_last;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last(9) <= PriceSummaryWriter_l_inst_l_count_order_bus_wdat_last;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data(BUS_DATA_WIDTH - 1 DOWNTO 0) <= PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_data;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data(BUS_DATA_WIDTH + BUS_DATA_WIDTH - 1 DOWNTO BUS_DATA_WIDTH) <= PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_data;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data(BUS_DATA_WIDTH * 2 + BUS_DATA_WIDTH - 1 DOWNTO BUS_DATA_WIDTH * 2) <= PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_data;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data(BUS_DATA_WIDTH * 3 + BUS_DATA_WIDTH - 1 DOWNTO BUS_DATA_WIDTH * 3) <= PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_data;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data(BUS_DATA_WIDTH * 4 + BUS_DATA_WIDTH - 1 DOWNTO BUS_DATA_WIDTH * 4) <= PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_data;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data(BUS_DATA_WIDTH * 5 + BUS_DATA_WIDTH - 1 DOWNTO BUS_DATA_WIDTH * 5) <= PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_data;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data(BUS_DATA_WIDTH * 6 + BUS_DATA_WIDTH - 1 DOWNTO BUS_DATA_WIDTH * 6) <= PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_data;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data(BUS_DATA_WIDTH * 7 + BUS_DATA_WIDTH - 1 DOWNTO BUS_DATA_WIDTH * 7) <= PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_data;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data(BUS_DATA_WIDTH * 8 + BUS_DATA_WIDTH - 1 DOWNTO BUS_DATA_WIDTH * 8) <= PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_data;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data(BUS_DATA_WIDTH * 9 + BUS_DATA_WIDTH - 1 DOWNTO BUS_DATA_WIDTH * 9) <= PriceSummaryWriter_l_inst_l_count_order_bus_wdat_data;
  PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_ready <= WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready(2);
  PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_ready <= WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready(2);
  PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_ready <= WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready(4);
  PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_ready <= WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready(4);
  PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_ready <= WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready(5);
  PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_ready <= WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready(5);
  PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_ready <= WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready(3);
  PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_ready <= WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready(3);
  PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_ready <= WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready(0);
  PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_ready <= WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready(0);
  PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_ready <= WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready(1);
  PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_ready <= WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready(1);
  PriceSummaryWriter_l_inst_l_count_order_bus_wreq_ready <= WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready(9);
  PriceSummaryWriter_l_inst_l_count_order_bus_wdat_ready <= WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready(9);
  PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_ready <= WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready(6);
  PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_ready <= WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready(6);
  PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_ready <= WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready(7);
  PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_ready <= WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready(7);
  PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_ready <= WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready(8);
  PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_ready <= WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready(8);
  RDAW64DW512LW8BS1BM16_inst : BusReadArbiterVec
  GENERIC MAP(
    BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
    BUS_DATA_WIDTH => BUS_DATA_WIDTH,
    BUS_LEN_WIDTH => BUS_LEN_WIDTH,
    NUM_SLAVE_PORTS => 7,
    ARB_METHOD => "RR-STICKY",
    MAX_OUTSTANDING => 4,
    RAM_CONFIG => "",
    SLV_REQ_SLICES => true,
    MST_REQ_SLICE => true,
    MST_DAT_SLICE => true,
    SLV_DAT_SLICES => true
  )
  PORT MAP(
    bcd_clk => bcd_clk,
    bcd_reset => bcd_reset,
    mst_rreq_valid => RDAW64DW512LW8BS1BM16_inst_mst_rreq_valid,
    mst_rreq_ready => RDAW64DW512LW8BS1BM16_inst_mst_rreq_ready,
    mst_rreq_addr => RDAW64DW512LW8BS1BM16_inst_mst_rreq_addr,
    mst_rreq_len => RDAW64DW512LW8BS1BM16_inst_mst_rreq_len,
    mst_rdat_valid => RDAW64DW512LW8BS1BM16_inst_mst_rdat_valid,
    mst_rdat_ready => RDAW64DW512LW8BS1BM16_inst_mst_rdat_ready,
    mst_rdat_data => RDAW64DW512LW8BS1BM16_inst_mst_rdat_data,
    mst_rdat_last => RDAW64DW512LW8BS1BM16_inst_mst_rdat_last,
    bsv_rreq_valid => RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid,
    bsv_rreq_ready => RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready,
    bsv_rreq_len => RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len,
    bsv_rreq_addr => RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr,
    bsv_rdat_valid => RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid,
    bsv_rdat_ready => RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready,
    bsv_rdat_last => RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last,
    bsv_rdat_data => RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data
  );

  rd_mst_rreq_valid <= RDAW64DW512LW8BS1BM16_inst_mst_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_mst_rreq_ready <= rd_mst_rreq_ready;
  rd_mst_rreq_addr <= RDAW64DW512LW8BS1BM16_inst_mst_rreq_addr;
  rd_mst_rreq_len <= RDAW64DW512LW8BS1BM16_inst_mst_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_mst_rdat_valid <= rd_mst_rdat_valid;
  rd_mst_rdat_ready <= RDAW64DW512LW8BS1BM16_inst_mst_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_mst_rdat_data <= rd_mst_rdat_data;
  RDAW64DW512LW8BS1BM16_inst_mst_rdat_last <= rd_mst_rdat_last;

  PriceSummary_Nucleus_inst_mmio_awvalid <= mmio_awvalid;
  mmio_awready <= PriceSummary_Nucleus_inst_mmio_awready;
  PriceSummary_Nucleus_inst_mmio_awaddr <= mmio_awaddr;
  PriceSummary_Nucleus_inst_mmio_wvalid <= mmio_wvalid;
  mmio_wready <= PriceSummary_Nucleus_inst_mmio_wready;
  PriceSummary_Nucleus_inst_mmio_wdata <= mmio_wdata;
  PriceSummary_Nucleus_inst_mmio_wstrb <= mmio_wstrb;
  mmio_bvalid <= PriceSummary_Nucleus_inst_mmio_bvalid;
  PriceSummary_Nucleus_inst_mmio_bready <= mmio_bready;
  mmio_bresp <= PriceSummary_Nucleus_inst_mmio_bresp;
  PriceSummary_Nucleus_inst_mmio_arvalid <= mmio_arvalid;
  mmio_arready <= PriceSummary_Nucleus_inst_mmio_arready;
  PriceSummary_Nucleus_inst_mmio_araddr <= mmio_araddr;
  mmio_rvalid <= PriceSummary_Nucleus_inst_mmio_rvalid;
  PriceSummary_Nucleus_inst_mmio_rready <= mmio_rready;
  mmio_rdata <= PriceSummary_Nucleus_inst_mmio_rdata;
  mmio_rresp <= PriceSummary_Nucleus_inst_mmio_rresp;

  PriceSummary_Nucleus_inst_l_quantity_valid <= PriceSummary_l_inst_l_quantity_valid;
  PriceSummary_l_inst_l_quantity_ready <= PriceSummary_Nucleus_inst_l_quantity_ready;
  PriceSummary_Nucleus_inst_l_quantity_dvalid <= PriceSummary_l_inst_l_quantity_dvalid;
  PriceSummary_Nucleus_inst_l_quantity_last <= PriceSummary_l_inst_l_quantity_last;
  PriceSummary_Nucleus_inst_l_quantity <= PriceSummary_l_inst_l_quantity;

  PriceSummary_Nucleus_inst_l_extendedprice_valid <= PriceSummary_l_inst_l_extendedprice_valid;
  PriceSummary_l_inst_l_extendedprice_ready <= PriceSummary_Nucleus_inst_l_extendedprice_ready;
  PriceSummary_Nucleus_inst_l_extendedprice_dvalid <= PriceSummary_l_inst_l_extendedprice_dvalid;
  PriceSummary_Nucleus_inst_l_extendedprice_last <= PriceSummary_l_inst_l_extendedprice_last;
  PriceSummary_Nucleus_inst_l_extendedprice <= PriceSummary_l_inst_l_extendedprice;

  PriceSummary_Nucleus_inst_l_discount_valid <= PriceSummary_l_inst_l_discount_valid;
  PriceSummary_l_inst_l_discount_ready <= PriceSummary_Nucleus_inst_l_discount_ready;
  PriceSummary_Nucleus_inst_l_discount_dvalid <= PriceSummary_l_inst_l_discount_dvalid;
  PriceSummary_Nucleus_inst_l_discount_last <= PriceSummary_l_inst_l_discount_last;
  PriceSummary_Nucleus_inst_l_discount <= PriceSummary_l_inst_l_discount;

  PriceSummary_Nucleus_inst_l_tax_valid <= PriceSummary_l_inst_l_tax_valid;
  PriceSummary_l_inst_l_tax_ready <= PriceSummary_Nucleus_inst_l_tax_ready;
  PriceSummary_Nucleus_inst_l_tax_dvalid <= PriceSummary_l_inst_l_tax_dvalid;
  PriceSummary_Nucleus_inst_l_tax_last <= PriceSummary_l_inst_l_tax_last;
  PriceSummary_Nucleus_inst_l_tax <= PriceSummary_l_inst_l_tax;

  PriceSummary_Nucleus_inst_l_returnflag_valid <= PriceSummary_l_inst_l_returnflag_valid;
  PriceSummary_l_inst_l_returnflag_ready <= PriceSummary_Nucleus_inst_l_returnflag_ready;
  PriceSummary_Nucleus_inst_l_returnflag_dvalid <= PriceSummary_l_inst_l_returnflag_dvalid;
  PriceSummary_Nucleus_inst_l_returnflag_last <= PriceSummary_l_inst_l_returnflag_last;
  PriceSummary_Nucleus_inst_l_returnflag_length <= PriceSummary_l_inst_l_returnflag_length;
  PriceSummary_Nucleus_inst_l_returnflag_count <= PriceSummary_l_inst_l_returnflag_count;
  PriceSummary_Nucleus_inst_l_returnflag_chars_valid <= PriceSummary_l_inst_l_returnflag_chars_valid;
  PriceSummary_l_inst_l_returnflag_chars_ready <= PriceSummary_Nucleus_inst_l_returnflag_chars_ready;
  PriceSummary_Nucleus_inst_l_returnflag_chars_dvalid <= PriceSummary_l_inst_l_returnflag_chars_dvalid;
  PriceSummary_Nucleus_inst_l_returnflag_chars_last <= PriceSummary_l_inst_l_returnflag_chars_last;
  PriceSummary_Nucleus_inst_l_returnflag_chars <= PriceSummary_l_inst_l_returnflag_chars;
  PriceSummary_Nucleus_inst_l_returnflag_chars_count <= PriceSummary_l_inst_l_returnflag_chars_count;

  PriceSummary_Nucleus_inst_l_linestatus_valid <= PriceSummary_l_inst_l_linestatus_valid;
  PriceSummary_l_inst_l_linestatus_ready <= PriceSummary_Nucleus_inst_l_linestatus_ready;
  PriceSummary_Nucleus_inst_l_linestatus_dvalid <= PriceSummary_l_inst_l_linestatus_dvalid;
  PriceSummary_Nucleus_inst_l_linestatus_last <= PriceSummary_l_inst_l_linestatus_last;
  PriceSummary_Nucleus_inst_l_linestatus_length <= PriceSummary_l_inst_l_linestatus_length;
  PriceSummary_Nucleus_inst_l_linestatus_count <= PriceSummary_l_inst_l_linestatus_count;
  PriceSummary_Nucleus_inst_l_linestatus_chars_valid <= PriceSummary_l_inst_l_linestatus_chars_valid;
  PriceSummary_l_inst_l_linestatus_chars_ready <= PriceSummary_Nucleus_inst_l_linestatus_chars_ready;
  PriceSummary_Nucleus_inst_l_linestatus_chars_dvalid <= PriceSummary_l_inst_l_linestatus_chars_dvalid;
  PriceSummary_Nucleus_inst_l_linestatus_chars_last <= PriceSummary_l_inst_l_linestatus_chars_last;
  PriceSummary_Nucleus_inst_l_linestatus_chars <= PriceSummary_l_inst_l_linestatus_chars;
  PriceSummary_Nucleus_inst_l_linestatus_chars_count <= PriceSummary_l_inst_l_linestatus_chars_count;

  PriceSummary_Nucleus_inst_l_shipdate_valid <= PriceSummary_l_inst_l_shipdate_valid;
  PriceSummary_l_inst_l_shipdate_ready <= PriceSummary_Nucleus_inst_l_shipdate_ready;
  PriceSummary_Nucleus_inst_l_shipdate_dvalid <= PriceSummary_l_inst_l_shipdate_dvalid;
  PriceSummary_Nucleus_inst_l_shipdate_last <= PriceSummary_l_inst_l_shipdate_last;
  PriceSummary_Nucleus_inst_l_shipdate <= PriceSummary_l_inst_l_shipdate;

  PriceSummary_Nucleus_inst_l_quantity_unl_valid <= PriceSummary_l_inst_l_quantity_unl_valid;
  PriceSummary_l_inst_l_quantity_unl_ready <= PriceSummary_Nucleus_inst_l_quantity_unl_ready;
  PriceSummary_Nucleus_inst_l_quantity_unl_tag <= PriceSummary_l_inst_l_quantity_unl_tag;

  PriceSummary_Nucleus_inst_l_extendedprice_unl_valid <= PriceSummary_l_inst_l_extendedprice_unl_valid;
  PriceSummary_l_inst_l_extendedprice_unl_ready <= PriceSummary_Nucleus_inst_l_extendedprice_unl_ready;
  PriceSummary_Nucleus_inst_l_extendedprice_unl_tag <= PriceSummary_l_inst_l_extendedprice_unl_tag;

  PriceSummary_Nucleus_inst_l_discount_unl_valid <= PriceSummary_l_inst_l_discount_unl_valid;
  PriceSummary_l_inst_l_discount_unl_ready <= PriceSummary_Nucleus_inst_l_discount_unl_ready;
  PriceSummary_Nucleus_inst_l_discount_unl_tag <= PriceSummary_l_inst_l_discount_unl_tag;

  PriceSummary_Nucleus_inst_l_tax_unl_valid <= PriceSummary_l_inst_l_tax_unl_valid;
  PriceSummary_l_inst_l_tax_unl_ready <= PriceSummary_Nucleus_inst_l_tax_unl_ready;
  PriceSummary_Nucleus_inst_l_tax_unl_tag <= PriceSummary_l_inst_l_tax_unl_tag;

  PriceSummary_Nucleus_inst_l_returnflag_unl_valid <= PriceSummary_l_inst_l_returnflag_unl_valid;
  PriceSummary_l_inst_l_returnflag_unl_ready <= PriceSummary_Nucleus_inst_l_returnflag_unl_ready;
  PriceSummary_Nucleus_inst_l_returnflag_unl_tag <= PriceSummary_l_inst_l_returnflag_unl_tag;

  PriceSummary_Nucleus_inst_l_linestatus_unl_valid <= PriceSummary_l_inst_l_linestatus_unl_valid;
  PriceSummary_l_inst_l_linestatus_unl_ready <= PriceSummary_Nucleus_inst_l_linestatus_unl_ready;
  PriceSummary_Nucleus_inst_l_linestatus_unl_tag <= PriceSummary_l_inst_l_linestatus_unl_tag;

  PriceSummary_Nucleus_inst_l_shipdate_unl_valid <= PriceSummary_l_inst_l_shipdate_unl_valid;
  PriceSummary_l_inst_l_shipdate_unl_ready <= PriceSummary_Nucleus_inst_l_shipdate_unl_ready;
  PriceSummary_Nucleus_inst_l_shipdate_unl_tag <= PriceSummary_l_inst_l_shipdate_unl_tag;

  PriceSummary_l_inst_l_quantity_cmd_valid <= PriceSummary_Nucleus_inst_l_quantity_cmd_valid;
  PriceSummary_Nucleus_inst_l_quantity_cmd_ready <= PriceSummary_l_inst_l_quantity_cmd_ready;
  PriceSummary_l_inst_l_quantity_cmd_firstIdx <= PriceSummary_Nucleus_inst_l_quantity_cmd_firstIdx;
  PriceSummary_l_inst_l_quantity_cmd_lastIdx <= PriceSummary_Nucleus_inst_l_quantity_cmd_lastIdx;
  PriceSummary_l_inst_l_quantity_cmd_ctrl <= PriceSummary_Nucleus_inst_l_quantity_cmd_ctrl;
  PriceSummary_l_inst_l_quantity_cmd_tag <= PriceSummary_Nucleus_inst_l_quantity_cmd_tag;

  PriceSummary_l_inst_l_extendedprice_cmd_valid <= PriceSummary_Nucleus_inst_l_extendedprice_cmd_valid;
  PriceSummary_Nucleus_inst_l_extendedprice_cmd_ready <= PriceSummary_l_inst_l_extendedprice_cmd_ready;
  PriceSummary_l_inst_l_extendedprice_cmd_firstIdx <= PriceSummary_Nucleus_inst_l_extendedprice_cmd_firstIdx;
  PriceSummary_l_inst_l_extendedprice_cmd_lastIdx <= PriceSummary_Nucleus_inst_l_extendedprice_cmd_lastIdx;
  PriceSummary_l_inst_l_extendedprice_cmd_ctrl <= PriceSummary_Nucleus_inst_l_extendedprice_cmd_ctrl;
  PriceSummary_l_inst_l_extendedprice_cmd_tag <= PriceSummary_Nucleus_inst_l_extendedprice_cmd_tag;

  PriceSummary_l_inst_l_discount_cmd_valid <= PriceSummary_Nucleus_inst_l_discount_cmd_valid;
  PriceSummary_Nucleus_inst_l_discount_cmd_ready <= PriceSummary_l_inst_l_discount_cmd_ready;
  PriceSummary_l_inst_l_discount_cmd_firstIdx <= PriceSummary_Nucleus_inst_l_discount_cmd_firstIdx;
  PriceSummary_l_inst_l_discount_cmd_lastIdx <= PriceSummary_Nucleus_inst_l_discount_cmd_lastIdx;
  PriceSummary_l_inst_l_discount_cmd_ctrl <= PriceSummary_Nucleus_inst_l_discount_cmd_ctrl;
  PriceSummary_l_inst_l_discount_cmd_tag <= PriceSummary_Nucleus_inst_l_discount_cmd_tag;

  PriceSummary_l_inst_l_tax_cmd_valid <= PriceSummary_Nucleus_inst_l_tax_cmd_valid;
  PriceSummary_Nucleus_inst_l_tax_cmd_ready <= PriceSummary_l_inst_l_tax_cmd_ready;
  PriceSummary_l_inst_l_tax_cmd_firstIdx <= PriceSummary_Nucleus_inst_l_tax_cmd_firstIdx;
  PriceSummary_l_inst_l_tax_cmd_lastIdx <= PriceSummary_Nucleus_inst_l_tax_cmd_lastIdx;
  PriceSummary_l_inst_l_tax_cmd_ctrl <= PriceSummary_Nucleus_inst_l_tax_cmd_ctrl;
  PriceSummary_l_inst_l_tax_cmd_tag <= PriceSummary_Nucleus_inst_l_tax_cmd_tag;

  PriceSummary_l_inst_l_returnflag_cmd_valid <= PriceSummary_Nucleus_inst_l_returnflag_cmd_valid;
  PriceSummary_Nucleus_inst_l_returnflag_cmd_ready <= PriceSummary_l_inst_l_returnflag_cmd_ready;
  PriceSummary_l_inst_l_returnflag_cmd_firstIdx <= PriceSummary_Nucleus_inst_l_returnflag_cmd_firstIdx;
  PriceSummary_l_inst_l_returnflag_cmd_lastIdx <= PriceSummary_Nucleus_inst_l_returnflag_cmd_lastIdx;
  PriceSummary_l_inst_l_returnflag_cmd_ctrl <= PriceSummary_Nucleus_inst_l_returnflag_cmd_ctrl;
  PriceSummary_l_inst_l_returnflag_cmd_tag <= PriceSummary_Nucleus_inst_l_returnflag_cmd_tag;

  PriceSummary_l_inst_l_linestatus_cmd_valid <= PriceSummary_Nucleus_inst_l_linestatus_cmd_valid;
  PriceSummary_Nucleus_inst_l_linestatus_cmd_ready <= PriceSummary_l_inst_l_linestatus_cmd_ready;
  PriceSummary_l_inst_l_linestatus_cmd_firstIdx <= PriceSummary_Nucleus_inst_l_linestatus_cmd_firstIdx;
  PriceSummary_l_inst_l_linestatus_cmd_lastIdx <= PriceSummary_Nucleus_inst_l_linestatus_cmd_lastIdx;
  PriceSummary_l_inst_l_linestatus_cmd_ctrl <= PriceSummary_Nucleus_inst_l_linestatus_cmd_ctrl;
  PriceSummary_l_inst_l_linestatus_cmd_tag <= PriceSummary_Nucleus_inst_l_linestatus_cmd_tag;

  PriceSummary_l_inst_l_shipdate_cmd_valid <= PriceSummary_Nucleus_inst_l_shipdate_cmd_valid;
  PriceSummary_Nucleus_inst_l_shipdate_cmd_ready <= PriceSummary_l_inst_l_shipdate_cmd_ready;
  PriceSummary_l_inst_l_shipdate_cmd_firstIdx <= PriceSummary_Nucleus_inst_l_shipdate_cmd_firstIdx;
  PriceSummary_l_inst_l_shipdate_cmd_lastIdx <= PriceSummary_Nucleus_inst_l_shipdate_cmd_lastIdx;
  PriceSummary_l_inst_l_shipdate_cmd_ctrl <= PriceSummary_Nucleus_inst_l_shipdate_cmd_ctrl;
  PriceSummary_l_inst_l_shipdate_cmd_tag <= PriceSummary_Nucleus_inst_l_shipdate_cmd_tag;

  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(0) <= PriceSummary_l_inst_l_quantity_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(1) <= PriceSummary_l_inst_l_extendedprice_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(2) <= PriceSummary_l_inst_l_discount_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(3) <= PriceSummary_l_inst_l_tax_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(4) <= PriceSummary_l_inst_l_returnflag_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(5) <= PriceSummary_l_inst_l_linestatus_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_valid(6) <= PriceSummary_l_inst_l_shipdate_bus_rreq_valid;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH - 1 DOWNTO 0) <= PriceSummary_l_inst_l_quantity_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH + BUS_LEN_WIDTH - 1 DOWNTO BUS_LEN_WIDTH) <= PriceSummary_l_inst_l_extendedprice_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH * 2 + BUS_LEN_WIDTH - 1 DOWNTO BUS_LEN_WIDTH * 2) <= PriceSummary_l_inst_l_discount_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH * 3 + BUS_LEN_WIDTH - 1 DOWNTO BUS_LEN_WIDTH * 3) <= PriceSummary_l_inst_l_tax_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH * 4 + BUS_LEN_WIDTH - 1 DOWNTO BUS_LEN_WIDTH * 4) <= PriceSummary_l_inst_l_returnflag_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH * 5 + BUS_LEN_WIDTH - 1 DOWNTO BUS_LEN_WIDTH * 5) <= PriceSummary_l_inst_l_linestatus_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_len(BUS_LEN_WIDTH * 6 + BUS_LEN_WIDTH - 1 DOWNTO BUS_LEN_WIDTH * 6) <= PriceSummary_l_inst_l_shipdate_bus_rreq_len;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH - 1 DOWNTO 0) <= PriceSummary_l_inst_l_quantity_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH + BUS_ADDR_WIDTH - 1 DOWNTO BUS_ADDR_WIDTH) <= PriceSummary_l_inst_l_extendedprice_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH * 2 + BUS_ADDR_WIDTH - 1 DOWNTO BUS_ADDR_WIDTH * 2) <= PriceSummary_l_inst_l_discount_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH * 3 + BUS_ADDR_WIDTH - 1 DOWNTO BUS_ADDR_WIDTH * 3) <= PriceSummary_l_inst_l_tax_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH * 4 + BUS_ADDR_WIDTH - 1 DOWNTO BUS_ADDR_WIDTH * 4) <= PriceSummary_l_inst_l_returnflag_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH * 5 + BUS_ADDR_WIDTH - 1 DOWNTO BUS_ADDR_WIDTH * 5) <= PriceSummary_l_inst_l_linestatus_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rreq_addr(BUS_ADDR_WIDTH * 6 + BUS_ADDR_WIDTH - 1 DOWNTO BUS_ADDR_WIDTH * 6) <= PriceSummary_l_inst_l_shipdate_bus_rreq_addr;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(0) <= PriceSummary_l_inst_l_quantity_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(1) <= PriceSummary_l_inst_l_extendedprice_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(2) <= PriceSummary_l_inst_l_discount_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(3) <= PriceSummary_l_inst_l_tax_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(4) <= PriceSummary_l_inst_l_returnflag_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(5) <= PriceSummary_l_inst_l_linestatus_bus_rdat_ready;
  RDAW64DW512LW8BS1BM16_inst_bsv_rdat_ready(6) <= PriceSummary_l_inst_l_shipdate_bus_rdat_ready;
  PriceSummary_l_inst_l_tax_bus_rreq_ready <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(3);
  PriceSummary_l_inst_l_tax_bus_rdat_valid <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(3);
  PriceSummary_l_inst_l_tax_bus_rdat_last <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(3);
  PriceSummary_l_inst_l_tax_bus_rdat_data <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH * 3 + BUS_DATA_WIDTH - 1 DOWNTO BUS_DATA_WIDTH * 3);
  PriceSummary_l_inst_l_shipdate_bus_rreq_ready <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(6);
  PriceSummary_l_inst_l_shipdate_bus_rdat_valid <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(6);
  PriceSummary_l_inst_l_shipdate_bus_rdat_last <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(6);
  PriceSummary_l_inst_l_shipdate_bus_rdat_data <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH * 6 + BUS_DATA_WIDTH - 1 DOWNTO BUS_DATA_WIDTH * 6);
  PriceSummary_l_inst_l_returnflag_bus_rreq_ready <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(4);
  PriceSummary_l_inst_l_returnflag_bus_rdat_valid <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(4);
  PriceSummary_l_inst_l_returnflag_bus_rdat_last <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(4);
  PriceSummary_l_inst_l_returnflag_bus_rdat_data <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH * 4 + BUS_DATA_WIDTH - 1 DOWNTO BUS_DATA_WIDTH * 4);
  PriceSummary_l_inst_l_quantity_bus_rreq_ready <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(0);
  PriceSummary_l_inst_l_quantity_bus_rdat_valid <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(0);
  PriceSummary_l_inst_l_quantity_bus_rdat_last <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(0);
  PriceSummary_l_inst_l_quantity_bus_rdat_data <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH - 1 DOWNTO 0);
  PriceSummary_l_inst_l_linestatus_bus_rreq_ready <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(5);
  PriceSummary_l_inst_l_linestatus_bus_rdat_valid <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(5);
  PriceSummary_l_inst_l_linestatus_bus_rdat_last <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(5);
  PriceSummary_l_inst_l_linestatus_bus_rdat_data <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH * 5 + BUS_DATA_WIDTH - 1 DOWNTO BUS_DATA_WIDTH * 5);
  PriceSummary_l_inst_l_extendedprice_bus_rreq_ready <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(1);
  PriceSummary_l_inst_l_extendedprice_bus_rdat_valid <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(1);
  PriceSummary_l_inst_l_extendedprice_bus_rdat_last <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(1);
  PriceSummary_l_inst_l_extendedprice_bus_rdat_data <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH + BUS_DATA_WIDTH - 1 DOWNTO BUS_DATA_WIDTH);
  PriceSummary_l_inst_l_discount_bus_rreq_ready <= RDAW64DW512LW8BS1BM16_inst_bsv_rreq_ready(2);
  PriceSummary_l_inst_l_discount_bus_rdat_valid <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_valid(2);
  PriceSummary_l_inst_l_discount_bus_rdat_last <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_last(2);
  PriceSummary_l_inst_l_discount_bus_rdat_data <= RDAW64DW512LW8BS1BM16_inst_bsv_rdat_data(BUS_DATA_WIDTH * 2 + BUS_DATA_WIDTH - 1 DOWNTO BUS_DATA_WIDTH * 2);

END ARCHITECTURE;