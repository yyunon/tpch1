-------------------------------------
-- Defines the dataPath width
--
-------------------------------------
package mypackage is
   constant XBITS :INTEGER := 64; 
   constant YBITS :INTEGER := 32;
   constant GRAIN :INTEGER := 4; --Number of add-sub cells
end mypackage;

