-- Copyright 2018-2019 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
-- This file was generated by Fletchgen. Modify this file at your own risk.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.Array_pkg.all;
use work.mmio_pkg.all;

entity PriceSummaryWriter_Nucleus is
  generic (
    INDEX_WIDTH                     : integer := 32;
    TAG_WIDTH                       : integer := 1;
    L_RETURNFLAG_O_BUS_ADDR_WIDTH   : integer := 64;
    L_LINESTATUS_O_BUS_ADDR_WIDTH   : integer := 64;
    L_SUM_QTY_BUS_ADDR_WIDTH        : integer := 64;
    L_SUM_BASE_PRICE_BUS_ADDR_WIDTH : integer := 64;
    L_SUM_DISC_PRICE_BUS_ADDR_WIDTH : integer := 64;
    L_SUM_CHARGE_BUS_ADDR_WIDTH     : integer := 64;
    L_AVG_QTY_BUS_ADDR_WIDTH        : integer := 64;
    L_AVG_PRICE_BUS_ADDR_WIDTH      : integer := 64;
    L_AVG_DISC_BUS_ADDR_WIDTH       : integer := 64;
    L_COUNT_ORDER_BUS_ADDR_WIDTH    : integer := 64
  );
  port (
    kcd_clk                       : in  std_logic;
    kcd_reset                     : in  std_logic;
    mmio_awvalid                  : in  std_logic;
    mmio_awready                  : out std_logic;
    mmio_awaddr                   : in  std_logic_vector(31 downto 0);
    mmio_wvalid                   : in  std_logic;
    mmio_wready                   : out std_logic;
    mmio_wdata                    : in  std_logic_vector(31 downto 0);
    mmio_wstrb                    : in  std_logic_vector(3 downto 0);
    mmio_bvalid                   : out std_logic;
    mmio_bready                   : in  std_logic;
    mmio_bresp                    : out std_logic_vector(1 downto 0);
    mmio_arvalid                  : in  std_logic;
    mmio_arready                  : out std_logic;
    mmio_araddr                   : in  std_logic_vector(31 downto 0);
    mmio_rvalid                   : out std_logic;
    mmio_rready                   : in  std_logic;
    mmio_rdata                    : out std_logic_vector(31 downto 0);
    mmio_rresp                    : out std_logic_vector(1 downto 0);
    l_returnflag_o_valid          : out std_logic;
    l_returnflag_o_ready          : in  std_logic;
    l_returnflag_o_dvalid         : out std_logic;
    l_returnflag_o_last           : out std_logic;
    l_returnflag_o_length         : out std_logic_vector(31 downto 0);
    l_returnflag_o_count          : out std_logic_vector(0 downto 0);
    l_returnflag_o_chars_valid    : out std_logic;
    l_returnflag_o_chars_ready    : in  std_logic;
    l_returnflag_o_chars_dvalid   : out std_logic;
    l_returnflag_o_chars_last     : out std_logic;
    l_returnflag_o_chars          : out std_logic_vector(7 downto 0);
    l_returnflag_o_chars_count    : out std_logic_vector(0 downto 0);
    l_linestatus_o_valid          : out std_logic;
    l_linestatus_o_ready          : in  std_logic;
    l_linestatus_o_dvalid         : out std_logic;
    l_linestatus_o_last           : out std_logic;
    l_linestatus_o_length         : out std_logic_vector(31 downto 0);
    l_linestatus_o_count          : out std_logic_vector(0 downto 0);
    l_linestatus_o_chars_valid    : out std_logic;
    l_linestatus_o_chars_ready    : in  std_logic;
    l_linestatus_o_chars_dvalid   : out std_logic;
    l_linestatus_o_chars_last     : out std_logic;
    l_linestatus_o_chars          : out std_logic_vector(7 downto 0);
    l_linestatus_o_chars_count    : out std_logic_vector(0 downto 0);
    l_sum_qty_valid               : out std_logic;
    l_sum_qty_ready               : in  std_logic;
    l_sum_qty_dvalid              : out std_logic;
    l_sum_qty_last                : out std_logic;
    l_sum_qty                     : out std_logic_vector(63 downto 0);
    l_sum_base_price_valid        : out std_logic;
    l_sum_base_price_ready        : in  std_logic;
    l_sum_base_price_dvalid       : out std_logic;
    l_sum_base_price_last         : out std_logic;
    l_sum_base_price              : out std_logic_vector(63 downto 0);
    l_sum_disc_price_valid        : out std_logic;
    l_sum_disc_price_ready        : in  std_logic;
    l_sum_disc_price_dvalid       : out std_logic;
    l_sum_disc_price_last         : out std_logic;
    l_sum_disc_price              : out std_logic_vector(63 downto 0);
    l_sum_charge_valid            : out std_logic;
    l_sum_charge_ready            : in  std_logic;
    l_sum_charge_dvalid           : out std_logic;
    l_sum_charge_last             : out std_logic;
    l_sum_charge                  : out std_logic_vector(63 downto 0);
    l_avg_qty_valid               : out std_logic;
    l_avg_qty_ready               : in  std_logic;
    l_avg_qty_dvalid              : out std_logic;
    l_avg_qty_last                : out std_logic;
    l_avg_qty                     : out std_logic_vector(63 downto 0);
    l_avg_price_valid             : out std_logic;
    l_avg_price_ready             : in  std_logic;
    l_avg_price_dvalid            : out std_logic;
    l_avg_price_last              : out std_logic;
    l_avg_price                   : out std_logic_vector(63 downto 0);
    l_avg_disc_valid              : out std_logic;
    l_avg_disc_ready              : in  std_logic;
    l_avg_disc_dvalid             : out std_logic;
    l_avg_disc_last               : out std_logic;
    l_avg_disc                    : out std_logic_vector(63 downto 0);
    l_count_order_valid           : out std_logic;
    l_count_order_ready           : in  std_logic;
    l_count_order_dvalid          : out std_logic;
    l_count_order_last            : out std_logic;
    l_count_order                 : out std_logic_vector(63 downto 0);
    l_returnflag_o_unl_valid      : in  std_logic;
    l_returnflag_o_unl_ready      : out std_logic;
    l_returnflag_o_unl_tag        : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_linestatus_o_unl_valid      : in  std_logic;
    l_linestatus_o_unl_ready      : out std_logic;
    l_linestatus_o_unl_tag        : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_sum_qty_unl_valid           : in  std_logic;
    l_sum_qty_unl_ready           : out std_logic;
    l_sum_qty_unl_tag             : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_sum_base_price_unl_valid    : in  std_logic;
    l_sum_base_price_unl_ready    : out std_logic;
    l_sum_base_price_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_sum_disc_price_unl_valid    : in  std_logic;
    l_sum_disc_price_unl_ready    : out std_logic;
    l_sum_disc_price_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_sum_charge_unl_valid        : in  std_logic;
    l_sum_charge_unl_ready        : out std_logic;
    l_sum_charge_unl_tag          : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_avg_qty_unl_valid           : in  std_logic;
    l_avg_qty_unl_ready           : out std_logic;
    l_avg_qty_unl_tag             : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_avg_price_unl_valid         : in  std_logic;
    l_avg_price_unl_ready         : out std_logic;
    l_avg_price_unl_tag           : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_avg_disc_unl_valid          : in  std_logic;
    l_avg_disc_unl_ready          : out std_logic;
    l_avg_disc_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_count_order_unl_valid       : in  std_logic;
    l_count_order_unl_ready       : out std_logic;
    l_count_order_unl_tag         : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_returnflag_o_cmd_valid      : out std_logic;
    l_returnflag_o_cmd_ready      : in  std_logic;
    l_returnflag_o_cmd_firstIdx   : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_returnflag_o_cmd_lastIdx    : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_returnflag_o_cmd_ctrl       : out std_logic_vector(L_RETURNFLAG_O_BUS_ADDR_WIDTH*2-1 downto 0);
    l_returnflag_o_cmd_tag        : out std_logic_vector(TAG_WIDTH-1 downto 0);
    l_linestatus_o_cmd_valid      : out std_logic;
    l_linestatus_o_cmd_ready      : in  std_logic;
    l_linestatus_o_cmd_firstIdx   : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_linestatus_o_cmd_lastIdx    : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_linestatus_o_cmd_ctrl       : out std_logic_vector(L_LINESTATUS_O_BUS_ADDR_WIDTH*2-1 downto 0);
    l_linestatus_o_cmd_tag        : out std_logic_vector(TAG_WIDTH-1 downto 0);
    l_sum_qty_cmd_valid           : out std_logic;
    l_sum_qty_cmd_ready           : in  std_logic;
    l_sum_qty_cmd_firstIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_sum_qty_cmd_lastIdx         : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_sum_qty_cmd_ctrl            : out std_logic_vector(L_SUM_QTY_BUS_ADDR_WIDTH-1 downto 0);
    l_sum_qty_cmd_tag             : out std_logic_vector(TAG_WIDTH-1 downto 0);
    l_sum_base_price_cmd_valid    : out std_logic;
    l_sum_base_price_cmd_ready    : in  std_logic;
    l_sum_base_price_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_sum_base_price_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_sum_base_price_cmd_ctrl     : out std_logic_vector(L_SUM_BASE_PRICE_BUS_ADDR_WIDTH-1 downto 0);
    l_sum_base_price_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
    l_sum_disc_price_cmd_valid    : out std_logic;
    l_sum_disc_price_cmd_ready    : in  std_logic;
    l_sum_disc_price_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_sum_disc_price_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_sum_disc_price_cmd_ctrl     : out std_logic_vector(L_SUM_DISC_PRICE_BUS_ADDR_WIDTH-1 downto 0);
    l_sum_disc_price_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
    l_sum_charge_cmd_valid        : out std_logic;
    l_sum_charge_cmd_ready        : in  std_logic;
    l_sum_charge_cmd_firstIdx     : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_sum_charge_cmd_lastIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_sum_charge_cmd_ctrl         : out std_logic_vector(L_SUM_CHARGE_BUS_ADDR_WIDTH-1 downto 0);
    l_sum_charge_cmd_tag          : out std_logic_vector(TAG_WIDTH-1 downto 0);
    l_avg_qty_cmd_valid           : out std_logic;
    l_avg_qty_cmd_ready           : in  std_logic;
    l_avg_qty_cmd_firstIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_avg_qty_cmd_lastIdx         : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_avg_qty_cmd_ctrl            : out std_logic_vector(L_AVG_QTY_BUS_ADDR_WIDTH-1 downto 0);
    l_avg_qty_cmd_tag             : out std_logic_vector(TAG_WIDTH-1 downto 0);
    l_avg_price_cmd_valid         : out std_logic;
    l_avg_price_cmd_ready         : in  std_logic;
    l_avg_price_cmd_firstIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_avg_price_cmd_lastIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_avg_price_cmd_ctrl          : out std_logic_vector(L_AVG_PRICE_BUS_ADDR_WIDTH-1 downto 0);
    l_avg_price_cmd_tag           : out std_logic_vector(TAG_WIDTH-1 downto 0);
    l_avg_disc_cmd_valid          : out std_logic;
    l_avg_disc_cmd_ready          : in  std_logic;
    l_avg_disc_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_avg_disc_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_avg_disc_cmd_ctrl           : out std_logic_vector(L_AVG_DISC_BUS_ADDR_WIDTH-1 downto 0);
    l_avg_disc_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
    l_count_order_cmd_valid       : out std_logic;
    l_count_order_cmd_ready       : in  std_logic;
    l_count_order_cmd_firstIdx    : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_count_order_cmd_lastIdx     : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_count_order_cmd_ctrl        : out std_logic_vector(L_COUNT_ORDER_BUS_ADDR_WIDTH-1 downto 0);
    l_count_order_cmd_tag         : out std_logic_vector(TAG_WIDTH-1 downto 0)
  );
end entity;

architecture Implementation of PriceSummaryWriter_Nucleus is
  component PriceSummaryWriter is
    generic (
      INDEX_WIDTH : integer := 32;
      TAG_WIDTH   : integer := 1
    );
    port (
      kcd_clk                       : in  std_logic;
      kcd_reset                     : in  std_logic;
      l_returnflag_o_valid          : out std_logic;
      l_returnflag_o_ready          : in  std_logic;
      l_returnflag_o_dvalid         : out std_logic;
      l_returnflag_o_last           : out std_logic;
      l_returnflag_o_length         : out std_logic_vector(31 downto 0);
      l_returnflag_o_count          : out std_logic_vector(0 downto 0);
      l_returnflag_o_chars_valid    : out std_logic;
      l_returnflag_o_chars_ready    : in  std_logic;
      l_returnflag_o_chars_dvalid   : out std_logic;
      l_returnflag_o_chars_last     : out std_logic;
      l_returnflag_o_chars          : out std_logic_vector(7 downto 0);
      l_returnflag_o_chars_count    : out std_logic_vector(0 downto 0);
      l_linestatus_o_valid          : out std_logic;
      l_linestatus_o_ready          : in  std_logic;
      l_linestatus_o_dvalid         : out std_logic;
      l_linestatus_o_last           : out std_logic;
      l_linestatus_o_length         : out std_logic_vector(31 downto 0);
      l_linestatus_o_count          : out std_logic_vector(0 downto 0);
      l_linestatus_o_chars_valid    : out std_logic;
      l_linestatus_o_chars_ready    : in  std_logic;
      l_linestatus_o_chars_dvalid   : out std_logic;
      l_linestatus_o_chars_last     : out std_logic;
      l_linestatus_o_chars          : out std_logic_vector(7 downto 0);
      l_linestatus_o_chars_count    : out std_logic_vector(0 downto 0);
      l_sum_qty_valid               : out std_logic;
      l_sum_qty_ready               : in  std_logic;
      l_sum_qty_dvalid              : out std_logic;
      l_sum_qty_last                : out std_logic;
      l_sum_qty                     : out std_logic_vector(63 downto 0);
      l_sum_base_price_valid        : out std_logic;
      l_sum_base_price_ready        : in  std_logic;
      l_sum_base_price_dvalid       : out std_logic;
      l_sum_base_price_last         : out std_logic;
      l_sum_base_price              : out std_logic_vector(63 downto 0);
      l_sum_disc_price_valid        : out std_logic;
      l_sum_disc_price_ready        : in  std_logic;
      l_sum_disc_price_dvalid       : out std_logic;
      l_sum_disc_price_last         : out std_logic;
      l_sum_disc_price              : out std_logic_vector(63 downto 0);
      l_sum_charge_valid            : out std_logic;
      l_sum_charge_ready            : in  std_logic;
      l_sum_charge_dvalid           : out std_logic;
      l_sum_charge_last             : out std_logic;
      l_sum_charge                  : out std_logic_vector(63 downto 0);
      l_avg_qty_valid               : out std_logic;
      l_avg_qty_ready               : in  std_logic;
      l_avg_qty_dvalid              : out std_logic;
      l_avg_qty_last                : out std_logic;
      l_avg_qty                     : out std_logic_vector(63 downto 0);
      l_avg_price_valid             : out std_logic;
      l_avg_price_ready             : in  std_logic;
      l_avg_price_dvalid            : out std_logic;
      l_avg_price_last              : out std_logic;
      l_avg_price                   : out std_logic_vector(63 downto 0);
      l_avg_disc_valid              : out std_logic;
      l_avg_disc_ready              : in  std_logic;
      l_avg_disc_dvalid             : out std_logic;
      l_avg_disc_last               : out std_logic;
      l_avg_disc                    : out std_logic_vector(63 downto 0);
      l_count_order_valid           : out std_logic;
      l_count_order_ready           : in  std_logic;
      l_count_order_dvalid          : out std_logic;
      l_count_order_last            : out std_logic;
      l_count_order                 : out std_logic_vector(63 downto 0);
      l_returnflag_o_unl_valid      : in  std_logic;
      l_returnflag_o_unl_ready      : out std_logic;
      l_returnflag_o_unl_tag        : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_linestatus_o_unl_valid      : in  std_logic;
      l_linestatus_o_unl_ready      : out std_logic;
      l_linestatus_o_unl_tag        : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_sum_qty_unl_valid           : in  std_logic;
      l_sum_qty_unl_ready           : out std_logic;
      l_sum_qty_unl_tag             : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_sum_base_price_unl_valid    : in  std_logic;
      l_sum_base_price_unl_ready    : out std_logic;
      l_sum_base_price_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_sum_disc_price_unl_valid    : in  std_logic;
      l_sum_disc_price_unl_ready    : out std_logic;
      l_sum_disc_price_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_sum_charge_unl_valid        : in  std_logic;
      l_sum_charge_unl_ready        : out std_logic;
      l_sum_charge_unl_tag          : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_avg_qty_unl_valid           : in  std_logic;
      l_avg_qty_unl_ready           : out std_logic;
      l_avg_qty_unl_tag             : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_avg_price_unl_valid         : in  std_logic;
      l_avg_price_unl_ready         : out std_logic;
      l_avg_price_unl_tag           : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_avg_disc_unl_valid          : in  std_logic;
      l_avg_disc_unl_ready          : out std_logic;
      l_avg_disc_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_count_order_unl_valid       : in  std_logic;
      l_count_order_unl_ready       : out std_logic;
      l_count_order_unl_tag         : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_returnflag_o_cmd_valid      : out std_logic;
      l_returnflag_o_cmd_ready      : in  std_logic;
      l_returnflag_o_cmd_firstIdx   : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_returnflag_o_cmd_lastIdx    : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_returnflag_o_cmd_tag        : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_linestatus_o_cmd_valid      : out std_logic;
      l_linestatus_o_cmd_ready      : in  std_logic;
      l_linestatus_o_cmd_firstIdx   : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_linestatus_o_cmd_lastIdx    : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_linestatus_o_cmd_tag        : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_sum_qty_cmd_valid           : out std_logic;
      l_sum_qty_cmd_ready           : in  std_logic;
      l_sum_qty_cmd_firstIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_sum_qty_cmd_lastIdx         : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_sum_qty_cmd_tag             : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_sum_base_price_cmd_valid    : out std_logic;
      l_sum_base_price_cmd_ready    : in  std_logic;
      l_sum_base_price_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_sum_base_price_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_sum_base_price_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_sum_disc_price_cmd_valid    : out std_logic;
      l_sum_disc_price_cmd_ready    : in  std_logic;
      l_sum_disc_price_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_sum_disc_price_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_sum_disc_price_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_sum_charge_cmd_valid        : out std_logic;
      l_sum_charge_cmd_ready        : in  std_logic;
      l_sum_charge_cmd_firstIdx     : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_sum_charge_cmd_lastIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_sum_charge_cmd_tag          : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_avg_qty_cmd_valid           : out std_logic;
      l_avg_qty_cmd_ready           : in  std_logic;
      l_avg_qty_cmd_firstIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_avg_qty_cmd_lastIdx         : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_avg_qty_cmd_tag             : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_avg_price_cmd_valid         : out std_logic;
      l_avg_price_cmd_ready         : in  std_logic;
      l_avg_price_cmd_firstIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_avg_price_cmd_lastIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_avg_price_cmd_tag           : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_avg_disc_cmd_valid          : out std_logic;
      l_avg_disc_cmd_ready          : in  std_logic;
      l_avg_disc_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_avg_disc_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_avg_disc_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_count_order_cmd_valid       : out std_logic;
      l_count_order_cmd_ready       : in  std_logic;
      l_count_order_cmd_firstIdx    : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_count_order_cmd_lastIdx     : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_count_order_cmd_tag         : out std_logic_vector(TAG_WIDTH-1 downto 0);
      start                         : in  std_logic;
      stop                          : in  std_logic;
      reset                         : in  std_logic;
      idle                          : out std_logic;
      busy                          : out std_logic;
      done                          : out std_logic;
      result                        : out std_logic_vector(63 downto 0);
      l_firstidx                    : in  std_logic_vector(31 downto 0);
      l_lastidx                     : in  std_logic_vector(31 downto 0)
    );
  end component;

  signal PriceSummaryWriter_inst_l_returnflag_o_valid          : std_logic;
  signal PriceSummaryWriter_inst_l_returnflag_o_ready          : std_logic;
  signal PriceSummaryWriter_inst_l_returnflag_o_dvalid         : std_logic;
  signal PriceSummaryWriter_inst_l_returnflag_o_last           : std_logic;
  signal PriceSummaryWriter_inst_l_returnflag_o_length         : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_inst_l_returnflag_o_count          : std_logic_vector(0 downto 0);
  signal PriceSummaryWriter_inst_l_returnflag_o_chars_valid    : std_logic;
  signal PriceSummaryWriter_inst_l_returnflag_o_chars_ready    : std_logic;
  signal PriceSummaryWriter_inst_l_returnflag_o_chars_dvalid   : std_logic;
  signal PriceSummaryWriter_inst_l_returnflag_o_chars_last     : std_logic;
  signal PriceSummaryWriter_inst_l_returnflag_o_chars          : std_logic_vector(7 downto 0);
  signal PriceSummaryWriter_inst_l_returnflag_o_chars_count    : std_logic_vector(0 downto 0);

  signal PriceSummaryWriter_inst_l_linestatus_o_valid          : std_logic;
  signal PriceSummaryWriter_inst_l_linestatus_o_ready          : std_logic;
  signal PriceSummaryWriter_inst_l_linestatus_o_dvalid         : std_logic;
  signal PriceSummaryWriter_inst_l_linestatus_o_last           : std_logic;
  signal PriceSummaryWriter_inst_l_linestatus_o_length         : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_inst_l_linestatus_o_count          : std_logic_vector(0 downto 0);
  signal PriceSummaryWriter_inst_l_linestatus_o_chars_valid    : std_logic;
  signal PriceSummaryWriter_inst_l_linestatus_o_chars_ready    : std_logic;
  signal PriceSummaryWriter_inst_l_linestatus_o_chars_dvalid   : std_logic;
  signal PriceSummaryWriter_inst_l_linestatus_o_chars_last     : std_logic;
  signal PriceSummaryWriter_inst_l_linestatus_o_chars          : std_logic_vector(7 downto 0);
  signal PriceSummaryWriter_inst_l_linestatus_o_chars_count    : std_logic_vector(0 downto 0);

  signal PriceSummaryWriter_inst_l_sum_qty_valid               : std_logic;
  signal PriceSummaryWriter_inst_l_sum_qty_ready               : std_logic;
  signal PriceSummaryWriter_inst_l_sum_qty_dvalid              : std_logic;
  signal PriceSummaryWriter_inst_l_sum_qty_last                : std_logic;
  signal PriceSummaryWriter_inst_l_sum_qty                     : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_inst_l_sum_base_price_valid        : std_logic;
  signal PriceSummaryWriter_inst_l_sum_base_price_ready        : std_logic;
  signal PriceSummaryWriter_inst_l_sum_base_price_dvalid       : std_logic;
  signal PriceSummaryWriter_inst_l_sum_base_price_last         : std_logic;
  signal PriceSummaryWriter_inst_l_sum_base_price              : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_inst_l_sum_disc_price_valid        : std_logic;
  signal PriceSummaryWriter_inst_l_sum_disc_price_ready        : std_logic;
  signal PriceSummaryWriter_inst_l_sum_disc_price_dvalid       : std_logic;
  signal PriceSummaryWriter_inst_l_sum_disc_price_last         : std_logic;
  signal PriceSummaryWriter_inst_l_sum_disc_price              : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_inst_l_sum_charge_valid            : std_logic;
  signal PriceSummaryWriter_inst_l_sum_charge_ready            : std_logic;
  signal PriceSummaryWriter_inst_l_sum_charge_dvalid           : std_logic;
  signal PriceSummaryWriter_inst_l_sum_charge_last             : std_logic;
  signal PriceSummaryWriter_inst_l_sum_charge                  : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_inst_l_avg_qty_valid               : std_logic;
  signal PriceSummaryWriter_inst_l_avg_qty_ready               : std_logic;
  signal PriceSummaryWriter_inst_l_avg_qty_dvalid              : std_logic;
  signal PriceSummaryWriter_inst_l_avg_qty_last                : std_logic;
  signal PriceSummaryWriter_inst_l_avg_qty                     : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_inst_l_avg_price_valid             : std_logic;
  signal PriceSummaryWriter_inst_l_avg_price_ready             : std_logic;
  signal PriceSummaryWriter_inst_l_avg_price_dvalid            : std_logic;
  signal PriceSummaryWriter_inst_l_avg_price_last              : std_logic;
  signal PriceSummaryWriter_inst_l_avg_price                   : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_inst_l_avg_disc_valid              : std_logic;
  signal PriceSummaryWriter_inst_l_avg_disc_ready              : std_logic;
  signal PriceSummaryWriter_inst_l_avg_disc_dvalid             : std_logic;
  signal PriceSummaryWriter_inst_l_avg_disc_last               : std_logic;
  signal PriceSummaryWriter_inst_l_avg_disc                    : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_inst_l_count_order_valid           : std_logic;
  signal PriceSummaryWriter_inst_l_count_order_ready           : std_logic;
  signal PriceSummaryWriter_inst_l_count_order_dvalid          : std_logic;
  signal PriceSummaryWriter_inst_l_count_order_last            : std_logic;
  signal PriceSummaryWriter_inst_l_count_order                 : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_inst_l_returnflag_o_unl_valid      : std_logic;
  signal PriceSummaryWriter_inst_l_returnflag_o_unl_ready      : std_logic;
  signal PriceSummaryWriter_inst_l_returnflag_o_unl_tag        : std_logic_vector(0 downto 0);

  signal PriceSummaryWriter_inst_l_linestatus_o_unl_valid      : std_logic;
  signal PriceSummaryWriter_inst_l_linestatus_o_unl_ready      : std_logic;
  signal PriceSummaryWriter_inst_l_linestatus_o_unl_tag        : std_logic_vector(0 downto 0);

  signal PriceSummaryWriter_inst_l_sum_qty_unl_valid           : std_logic;
  signal PriceSummaryWriter_inst_l_sum_qty_unl_ready           : std_logic;
  signal PriceSummaryWriter_inst_l_sum_qty_unl_tag             : std_logic_vector(0 downto 0);

  signal PriceSummaryWriter_inst_l_sum_base_price_unl_valid    : std_logic;
  signal PriceSummaryWriter_inst_l_sum_base_price_unl_ready    : std_logic;
  signal PriceSummaryWriter_inst_l_sum_base_price_unl_tag      : std_logic_vector(0 downto 0);

  signal PriceSummaryWriter_inst_l_sum_disc_price_unl_valid    : std_logic;
  signal PriceSummaryWriter_inst_l_sum_disc_price_unl_ready    : std_logic;
  signal PriceSummaryWriter_inst_l_sum_disc_price_unl_tag      : std_logic_vector(0 downto 0);

  signal PriceSummaryWriter_inst_l_sum_charge_unl_valid        : std_logic;
  signal PriceSummaryWriter_inst_l_sum_charge_unl_ready        : std_logic;
  signal PriceSummaryWriter_inst_l_sum_charge_unl_tag          : std_logic_vector(0 downto 0);

  signal PriceSummaryWriter_inst_l_avg_qty_unl_valid           : std_logic;
  signal PriceSummaryWriter_inst_l_avg_qty_unl_ready           : std_logic;
  signal PriceSummaryWriter_inst_l_avg_qty_unl_tag             : std_logic_vector(0 downto 0);

  signal PriceSummaryWriter_inst_l_avg_price_unl_valid         : std_logic;
  signal PriceSummaryWriter_inst_l_avg_price_unl_ready         : std_logic;
  signal PriceSummaryWriter_inst_l_avg_price_unl_tag           : std_logic_vector(0 downto 0);

  signal PriceSummaryWriter_inst_l_avg_disc_unl_valid          : std_logic;
  signal PriceSummaryWriter_inst_l_avg_disc_unl_ready          : std_logic;
  signal PriceSummaryWriter_inst_l_avg_disc_unl_tag            : std_logic_vector(0 downto 0);

  signal PriceSummaryWriter_inst_l_count_order_unl_valid       : std_logic;
  signal PriceSummaryWriter_inst_l_count_order_unl_ready       : std_logic;
  signal PriceSummaryWriter_inst_l_count_order_unl_tag         : std_logic_vector(0 downto 0);

  signal PriceSummaryWriter_inst_l_returnflag_o_cmd_valid      : std_logic;
  signal PriceSummaryWriter_inst_l_returnflag_o_cmd_ready      : std_logic;
  signal PriceSummaryWriter_inst_l_returnflag_o_cmd_firstIdx   : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_inst_l_returnflag_o_cmd_lastIdx    : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_inst_l_returnflag_o_cmd_tag        : std_logic_vector(0 downto 0);

  signal PriceSummaryWriter_inst_l_linestatus_o_cmd_valid      : std_logic;
  signal PriceSummaryWriter_inst_l_linestatus_o_cmd_ready      : std_logic;
  signal PriceSummaryWriter_inst_l_linestatus_o_cmd_firstIdx   : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_inst_l_linestatus_o_cmd_lastIdx    : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_inst_l_linestatus_o_cmd_tag        : std_logic_vector(0 downto 0);

  signal PriceSummaryWriter_inst_l_sum_qty_cmd_valid           : std_logic;
  signal PriceSummaryWriter_inst_l_sum_qty_cmd_ready           : std_logic;
  signal PriceSummaryWriter_inst_l_sum_qty_cmd_firstIdx        : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_inst_l_sum_qty_cmd_lastIdx         : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_inst_l_sum_qty_cmd_tag             : std_logic_vector(0 downto 0);

  signal PriceSummaryWriter_inst_l_sum_base_price_cmd_valid    : std_logic;
  signal PriceSummaryWriter_inst_l_sum_base_price_cmd_ready    : std_logic;
  signal PriceSummaryWriter_inst_l_sum_base_price_cmd_firstIdx : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_inst_l_sum_base_price_cmd_lastIdx  : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_inst_l_sum_base_price_cmd_tag      : std_logic_vector(0 downto 0);

  signal PriceSummaryWriter_inst_l_sum_disc_price_cmd_valid    : std_logic;
  signal PriceSummaryWriter_inst_l_sum_disc_price_cmd_ready    : std_logic;
  signal PriceSummaryWriter_inst_l_sum_disc_price_cmd_firstIdx : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_inst_l_sum_disc_price_cmd_lastIdx  : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_inst_l_sum_disc_price_cmd_tag      : std_logic_vector(0 downto 0);

  signal PriceSummaryWriter_inst_l_sum_charge_cmd_valid        : std_logic;
  signal PriceSummaryWriter_inst_l_sum_charge_cmd_ready        : std_logic;
  signal PriceSummaryWriter_inst_l_sum_charge_cmd_firstIdx     : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_inst_l_sum_charge_cmd_lastIdx      : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_inst_l_sum_charge_cmd_tag          : std_logic_vector(0 downto 0);

  signal PriceSummaryWriter_inst_l_avg_qty_cmd_valid           : std_logic;
  signal PriceSummaryWriter_inst_l_avg_qty_cmd_ready           : std_logic;
  signal PriceSummaryWriter_inst_l_avg_qty_cmd_firstIdx        : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_inst_l_avg_qty_cmd_lastIdx         : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_inst_l_avg_qty_cmd_tag             : std_logic_vector(0 downto 0);

  signal PriceSummaryWriter_inst_l_avg_price_cmd_valid         : std_logic;
  signal PriceSummaryWriter_inst_l_avg_price_cmd_ready         : std_logic;
  signal PriceSummaryWriter_inst_l_avg_price_cmd_firstIdx      : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_inst_l_avg_price_cmd_lastIdx       : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_inst_l_avg_price_cmd_tag           : std_logic_vector(0 downto 0);

  signal PriceSummaryWriter_inst_l_avg_disc_cmd_valid          : std_logic;
  signal PriceSummaryWriter_inst_l_avg_disc_cmd_ready          : std_logic;
  signal PriceSummaryWriter_inst_l_avg_disc_cmd_firstIdx       : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_inst_l_avg_disc_cmd_lastIdx        : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_inst_l_avg_disc_cmd_tag            : std_logic_vector(0 downto 0);

  signal PriceSummaryWriter_inst_l_count_order_cmd_valid       : std_logic;
  signal PriceSummaryWriter_inst_l_count_order_cmd_ready       : std_logic;
  signal PriceSummaryWriter_inst_l_count_order_cmd_firstIdx    : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_inst_l_count_order_cmd_lastIdx     : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_inst_l_count_order_cmd_tag         : std_logic_vector(0 downto 0);

  signal PriceSummaryWriter_inst_start                         : std_logic;
  signal PriceSummaryWriter_inst_stop                          : std_logic;
  signal PriceSummaryWriter_inst_reset                         : std_logic;
  signal PriceSummaryWriter_inst_idle                          : std_logic;
  signal PriceSummaryWriter_inst_busy                          : std_logic;
  signal PriceSummaryWriter_inst_done                          : std_logic;
  signal PriceSummaryWriter_inst_result                        : std_logic_vector(63 downto 0);
  signal PriceSummaryWriter_inst_l_firstidx                    : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_inst_l_lastidx                     : std_logic_vector(31 downto 0);
  signal mmio_inst_f_start_data                                : std_logic;
  signal mmio_inst_f_stop_data                                 : std_logic;
  signal mmio_inst_f_reset_data                                : std_logic;
  signal mmio_inst_f_idle_write_data                           : std_logic;
  signal mmio_inst_f_busy_write_data                           : std_logic;
  signal mmio_inst_f_done_write_data                           : std_logic;
  signal mmio_inst_f_result_write_data                         : std_logic_vector(63 downto 0);
  signal mmio_inst_f_l_firstidx_data                           : std_logic_vector(31 downto 0);
  signal mmio_inst_f_l_lastidx_data                            : std_logic_vector(31 downto 0);
  signal mmio_inst_f_l_returnflag_o_offsets_data               : std_logic_vector(63 downto 0);
  signal mmio_inst_f_l_returnflag_o_values_data                : std_logic_vector(63 downto 0);
  signal mmio_inst_f_l_linestatus_o_offsets_data               : std_logic_vector(63 downto 0);
  signal mmio_inst_f_l_linestatus_o_values_data                : std_logic_vector(63 downto 0);
  signal mmio_inst_f_l_sum_qty_values_data                     : std_logic_vector(63 downto 0);
  signal mmio_inst_f_l_sum_base_price_values_data              : std_logic_vector(63 downto 0);
  signal mmio_inst_f_l_sum_disc_price_values_data              : std_logic_vector(63 downto 0);
  signal mmio_inst_f_l_sum_charge_values_data                  : std_logic_vector(63 downto 0);
  signal mmio_inst_f_l_avg_qty_values_data                     : std_logic_vector(63 downto 0);
  signal mmio_inst_f_l_avg_price_values_data                   : std_logic_vector(63 downto 0);
  signal mmio_inst_f_l_avg_disc_values_data                    : std_logic_vector(63 downto 0);
  signal mmio_inst_f_l_count_order_values_data                 : std_logic_vector(63 downto 0);
  signal mmio_inst_f_Profile_enable_data                       : std_logic;
  signal mmio_inst_f_Profile_clear_data                        : std_logic;
  signal mmio_inst_mmio_awvalid                                : std_logic;
  signal mmio_inst_mmio_awready                                : std_logic;
  signal mmio_inst_mmio_awaddr                                 : std_logic_vector(31 downto 0);
  signal mmio_inst_mmio_wvalid                                 : std_logic;
  signal mmio_inst_mmio_wready                                 : std_logic;
  signal mmio_inst_mmio_wdata                                  : std_logic_vector(31 downto 0);
  signal mmio_inst_mmio_wstrb                                  : std_logic_vector(3 downto 0);
  signal mmio_inst_mmio_bvalid                                 : std_logic;
  signal mmio_inst_mmio_bready                                 : std_logic;
  signal mmio_inst_mmio_bresp                                  : std_logic_vector(1 downto 0);
  signal mmio_inst_mmio_arvalid                                : std_logic;
  signal mmio_inst_mmio_arready                                : std_logic;
  signal mmio_inst_mmio_araddr                                 : std_logic_vector(31 downto 0);
  signal mmio_inst_mmio_rvalid                                 : std_logic;
  signal mmio_inst_mmio_rready                                 : std_logic;
  signal mmio_inst_mmio_rdata                                  : std_logic_vector(31 downto 0);
  signal mmio_inst_mmio_rresp                                  : std_logic_vector(1 downto 0);

  signal l_returnflag_o_cmd_accm_inst_kernel_cmd_valid         : std_logic;
  signal l_returnflag_o_cmd_accm_inst_kernel_cmd_ready         : std_logic;
  signal l_returnflag_o_cmd_accm_inst_kernel_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_returnflag_o_cmd_accm_inst_kernel_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_returnflag_o_cmd_accm_inst_kernel_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_returnflag_o_cmd_accm_inst_nucleus_cmd_valid        : std_logic;
  signal l_returnflag_o_cmd_accm_inst_nucleus_cmd_ready        : std_logic;
  signal l_returnflag_o_cmd_accm_inst_nucleus_cmd_firstIdx     : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_returnflag_o_cmd_accm_inst_nucleus_cmd_lastIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_returnflag_o_cmd_accm_inst_nucleus_cmd_ctrl         : std_logic_vector(2*L_RETURNFLAG_O_BUS_ADDR_WIDTH-1 downto 0);
  signal l_returnflag_o_cmd_accm_inst_nucleus_cmd_tag          : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_linestatus_o_cmd_accm_inst_kernel_cmd_valid         : std_logic;
  signal l_linestatus_o_cmd_accm_inst_kernel_cmd_ready         : std_logic;
  signal l_linestatus_o_cmd_accm_inst_kernel_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_linestatus_o_cmd_accm_inst_kernel_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_linestatus_o_cmd_accm_inst_kernel_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_linestatus_o_cmd_accm_inst_nucleus_cmd_valid        : std_logic;
  signal l_linestatus_o_cmd_accm_inst_nucleus_cmd_ready        : std_logic;
  signal l_linestatus_o_cmd_accm_inst_nucleus_cmd_firstIdx     : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_linestatus_o_cmd_accm_inst_nucleus_cmd_lastIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_linestatus_o_cmd_accm_inst_nucleus_cmd_ctrl         : std_logic_vector(2*L_LINESTATUS_O_BUS_ADDR_WIDTH-1 downto 0);
  signal l_linestatus_o_cmd_accm_inst_nucleus_cmd_tag          : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_sum_qty_cmd_accm_inst_kernel_cmd_valid              : std_logic;
  signal l_sum_qty_cmd_accm_inst_kernel_cmd_ready              : std_logic;
  signal l_sum_qty_cmd_accm_inst_kernel_cmd_firstIdx           : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_sum_qty_cmd_accm_inst_kernel_cmd_lastIdx            : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_sum_qty_cmd_accm_inst_kernel_cmd_tag                : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_sum_qty_cmd_accm_inst_nucleus_cmd_valid             : std_logic;
  signal l_sum_qty_cmd_accm_inst_nucleus_cmd_ready             : std_logic;
  signal l_sum_qty_cmd_accm_inst_nucleus_cmd_firstIdx          : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_sum_qty_cmd_accm_inst_nucleus_cmd_lastIdx           : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_sum_qty_cmd_accm_inst_nucleus_cmd_ctrl              : std_logic_vector(L_SUM_QTY_BUS_ADDR_WIDTH-1 downto 0);
  signal l_sum_qty_cmd_accm_inst_nucleus_cmd_tag               : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_sum_base_price_cmd_accm_inst_kernel_cmd_valid       : std_logic;
  signal l_sum_base_price_cmd_accm_inst_kernel_cmd_ready       : std_logic;
  signal l_sum_base_price_cmd_accm_inst_kernel_cmd_firstIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_sum_base_price_cmd_accm_inst_kernel_cmd_lastIdx     : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_sum_base_price_cmd_accm_inst_kernel_cmd_tag         : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_sum_base_price_cmd_accm_inst_nucleus_cmd_valid      : std_logic;
  signal l_sum_base_price_cmd_accm_inst_nucleus_cmd_ready      : std_logic;
  signal l_sum_base_price_cmd_accm_inst_nucleus_cmd_firstIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_sum_base_price_cmd_accm_inst_nucleus_cmd_lastIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_sum_base_price_cmd_accm_inst_nucleus_cmd_ctrl       : std_logic_vector(L_SUM_BASE_PRICE_BUS_ADDR_WIDTH-1 downto 0);
  signal l_sum_base_price_cmd_accm_inst_nucleus_cmd_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_sum_disc_price_cmd_accm_inst_kernel_cmd_valid       : std_logic;
  signal l_sum_disc_price_cmd_accm_inst_kernel_cmd_ready       : std_logic;
  signal l_sum_disc_price_cmd_accm_inst_kernel_cmd_firstIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_sum_disc_price_cmd_accm_inst_kernel_cmd_lastIdx     : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_sum_disc_price_cmd_accm_inst_kernel_cmd_tag         : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_sum_disc_price_cmd_accm_inst_nucleus_cmd_valid      : std_logic;
  signal l_sum_disc_price_cmd_accm_inst_nucleus_cmd_ready      : std_logic;
  signal l_sum_disc_price_cmd_accm_inst_nucleus_cmd_firstIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_sum_disc_price_cmd_accm_inst_nucleus_cmd_lastIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_sum_disc_price_cmd_accm_inst_nucleus_cmd_ctrl       : std_logic_vector(L_SUM_DISC_PRICE_BUS_ADDR_WIDTH-1 downto 0);
  signal l_sum_disc_price_cmd_accm_inst_nucleus_cmd_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_sum_charge_cmd_accm_inst_kernel_cmd_valid           : std_logic;
  signal l_sum_charge_cmd_accm_inst_kernel_cmd_ready           : std_logic;
  signal l_sum_charge_cmd_accm_inst_kernel_cmd_firstIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_sum_charge_cmd_accm_inst_kernel_cmd_lastIdx         : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_sum_charge_cmd_accm_inst_kernel_cmd_tag             : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_sum_charge_cmd_accm_inst_nucleus_cmd_valid          : std_logic;
  signal l_sum_charge_cmd_accm_inst_nucleus_cmd_ready          : std_logic;
  signal l_sum_charge_cmd_accm_inst_nucleus_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_sum_charge_cmd_accm_inst_nucleus_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_sum_charge_cmd_accm_inst_nucleus_cmd_ctrl           : std_logic_vector(L_SUM_CHARGE_BUS_ADDR_WIDTH-1 downto 0);
  signal l_sum_charge_cmd_accm_inst_nucleus_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_avg_qty_cmd_accm_inst_kernel_cmd_valid              : std_logic;
  signal l_avg_qty_cmd_accm_inst_kernel_cmd_ready              : std_logic;
  signal l_avg_qty_cmd_accm_inst_kernel_cmd_firstIdx           : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_avg_qty_cmd_accm_inst_kernel_cmd_lastIdx            : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_avg_qty_cmd_accm_inst_kernel_cmd_tag                : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_avg_qty_cmd_accm_inst_nucleus_cmd_valid             : std_logic;
  signal l_avg_qty_cmd_accm_inst_nucleus_cmd_ready             : std_logic;
  signal l_avg_qty_cmd_accm_inst_nucleus_cmd_firstIdx          : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_avg_qty_cmd_accm_inst_nucleus_cmd_lastIdx           : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_avg_qty_cmd_accm_inst_nucleus_cmd_ctrl              : std_logic_vector(L_AVG_QTY_BUS_ADDR_WIDTH-1 downto 0);
  signal l_avg_qty_cmd_accm_inst_nucleus_cmd_tag               : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_avg_price_cmd_accm_inst_kernel_cmd_valid            : std_logic;
  signal l_avg_price_cmd_accm_inst_kernel_cmd_ready            : std_logic;
  signal l_avg_price_cmd_accm_inst_kernel_cmd_firstIdx         : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_avg_price_cmd_accm_inst_kernel_cmd_lastIdx          : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_avg_price_cmd_accm_inst_kernel_cmd_tag              : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_avg_price_cmd_accm_inst_nucleus_cmd_valid           : std_logic;
  signal l_avg_price_cmd_accm_inst_nucleus_cmd_ready           : std_logic;
  signal l_avg_price_cmd_accm_inst_nucleus_cmd_firstIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_avg_price_cmd_accm_inst_nucleus_cmd_lastIdx         : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_avg_price_cmd_accm_inst_nucleus_cmd_ctrl            : std_logic_vector(L_AVG_PRICE_BUS_ADDR_WIDTH-1 downto 0);
  signal l_avg_price_cmd_accm_inst_nucleus_cmd_tag             : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_avg_disc_cmd_accm_inst_kernel_cmd_valid             : std_logic;
  signal l_avg_disc_cmd_accm_inst_kernel_cmd_ready             : std_logic;
  signal l_avg_disc_cmd_accm_inst_kernel_cmd_firstIdx          : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_avg_disc_cmd_accm_inst_kernel_cmd_lastIdx           : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_avg_disc_cmd_accm_inst_kernel_cmd_tag               : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_avg_disc_cmd_accm_inst_nucleus_cmd_valid            : std_logic;
  signal l_avg_disc_cmd_accm_inst_nucleus_cmd_ready            : std_logic;
  signal l_avg_disc_cmd_accm_inst_nucleus_cmd_firstIdx         : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_avg_disc_cmd_accm_inst_nucleus_cmd_lastIdx          : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_avg_disc_cmd_accm_inst_nucleus_cmd_ctrl             : std_logic_vector(L_AVG_DISC_BUS_ADDR_WIDTH-1 downto 0);
  signal l_avg_disc_cmd_accm_inst_nucleus_cmd_tag              : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_count_order_cmd_accm_inst_kernel_cmd_valid          : std_logic;
  signal l_count_order_cmd_accm_inst_kernel_cmd_ready          : std_logic;
  signal l_count_order_cmd_accm_inst_kernel_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_count_order_cmd_accm_inst_kernel_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_count_order_cmd_accm_inst_kernel_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_count_order_cmd_accm_inst_nucleus_cmd_valid         : std_logic;
  signal l_count_order_cmd_accm_inst_nucleus_cmd_ready         : std_logic;
  signal l_count_order_cmd_accm_inst_nucleus_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_count_order_cmd_accm_inst_nucleus_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_count_order_cmd_accm_inst_nucleus_cmd_ctrl          : std_logic_vector(L_COUNT_ORDER_BUS_ADDR_WIDTH-1 downto 0);
  signal l_count_order_cmd_accm_inst_nucleus_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_returnflag_o_cmd_accm_inst_ctrl   : std_logic_vector(2*L_RETURNFLAG_O_BUS_ADDR_WIDTH-1 downto 0);
  signal l_linestatus_o_cmd_accm_inst_ctrl   : std_logic_vector(2*L_LINESTATUS_O_BUS_ADDR_WIDTH-1 downto 0);
  signal l_sum_qty_cmd_accm_inst_ctrl        : std_logic_vector(L_SUM_QTY_BUS_ADDR_WIDTH-1 downto 0);
  signal l_sum_base_price_cmd_accm_inst_ctrl : std_logic_vector(L_SUM_BASE_PRICE_BUS_ADDR_WIDTH-1 downto 0);
  signal l_sum_disc_price_cmd_accm_inst_ctrl : std_logic_vector(L_SUM_DISC_PRICE_BUS_ADDR_WIDTH-1 downto 0);
  signal l_sum_charge_cmd_accm_inst_ctrl     : std_logic_vector(L_SUM_CHARGE_BUS_ADDR_WIDTH-1 downto 0);
  signal l_avg_qty_cmd_accm_inst_ctrl        : std_logic_vector(L_AVG_QTY_BUS_ADDR_WIDTH-1 downto 0);
  signal l_avg_price_cmd_accm_inst_ctrl      : std_logic_vector(L_AVG_PRICE_BUS_ADDR_WIDTH-1 downto 0);
  signal l_avg_disc_cmd_accm_inst_ctrl       : std_logic_vector(L_AVG_DISC_BUS_ADDR_WIDTH-1 downto 0);
  signal l_count_order_cmd_accm_inst_ctrl    : std_logic_vector(L_COUNT_ORDER_BUS_ADDR_WIDTH-1 downto 0);

begin
  PriceSummaryWriter_inst : PriceSummaryWriter
    generic map (
      INDEX_WIDTH => 32,
      TAG_WIDTH   => 1
    )
    port map (
      kcd_clk                       => kcd_clk,
      kcd_reset                     => kcd_reset,
      l_returnflag_o_valid          => PriceSummaryWriter_inst_l_returnflag_o_valid,
      l_returnflag_o_ready          => PriceSummaryWriter_inst_l_returnflag_o_ready,
      l_returnflag_o_dvalid         => PriceSummaryWriter_inst_l_returnflag_o_dvalid,
      l_returnflag_o_last           => PriceSummaryWriter_inst_l_returnflag_o_last,
      l_returnflag_o_length         => PriceSummaryWriter_inst_l_returnflag_o_length,
      l_returnflag_o_count          => PriceSummaryWriter_inst_l_returnflag_o_count,
      l_returnflag_o_chars_valid    => PriceSummaryWriter_inst_l_returnflag_o_chars_valid,
      l_returnflag_o_chars_ready    => PriceSummaryWriter_inst_l_returnflag_o_chars_ready,
      l_returnflag_o_chars_dvalid   => PriceSummaryWriter_inst_l_returnflag_o_chars_dvalid,
      l_returnflag_o_chars_last     => PriceSummaryWriter_inst_l_returnflag_o_chars_last,
      l_returnflag_o_chars          => PriceSummaryWriter_inst_l_returnflag_o_chars,
      l_returnflag_o_chars_count    => PriceSummaryWriter_inst_l_returnflag_o_chars_count,
      l_linestatus_o_valid          => PriceSummaryWriter_inst_l_linestatus_o_valid,
      l_linestatus_o_ready          => PriceSummaryWriter_inst_l_linestatus_o_ready,
      l_linestatus_o_dvalid         => PriceSummaryWriter_inst_l_linestatus_o_dvalid,
      l_linestatus_o_last           => PriceSummaryWriter_inst_l_linestatus_o_last,
      l_linestatus_o_length         => PriceSummaryWriter_inst_l_linestatus_o_length,
      l_linestatus_o_count          => PriceSummaryWriter_inst_l_linestatus_o_count,
      l_linestatus_o_chars_valid    => PriceSummaryWriter_inst_l_linestatus_o_chars_valid,
      l_linestatus_o_chars_ready    => PriceSummaryWriter_inst_l_linestatus_o_chars_ready,
      l_linestatus_o_chars_dvalid   => PriceSummaryWriter_inst_l_linestatus_o_chars_dvalid,
      l_linestatus_o_chars_last     => PriceSummaryWriter_inst_l_linestatus_o_chars_last,
      l_linestatus_o_chars          => PriceSummaryWriter_inst_l_linestatus_o_chars,
      l_linestatus_o_chars_count    => PriceSummaryWriter_inst_l_linestatus_o_chars_count,
      l_sum_qty_valid               => PriceSummaryWriter_inst_l_sum_qty_valid,
      l_sum_qty_ready               => PriceSummaryWriter_inst_l_sum_qty_ready,
      l_sum_qty_dvalid              => PriceSummaryWriter_inst_l_sum_qty_dvalid,
      l_sum_qty_last                => PriceSummaryWriter_inst_l_sum_qty_last,
      l_sum_qty                     => PriceSummaryWriter_inst_l_sum_qty,
      l_sum_base_price_valid        => PriceSummaryWriter_inst_l_sum_base_price_valid,
      l_sum_base_price_ready        => PriceSummaryWriter_inst_l_sum_base_price_ready,
      l_sum_base_price_dvalid       => PriceSummaryWriter_inst_l_sum_base_price_dvalid,
      l_sum_base_price_last         => PriceSummaryWriter_inst_l_sum_base_price_last,
      l_sum_base_price              => PriceSummaryWriter_inst_l_sum_base_price,
      l_sum_disc_price_valid        => PriceSummaryWriter_inst_l_sum_disc_price_valid,
      l_sum_disc_price_ready        => PriceSummaryWriter_inst_l_sum_disc_price_ready,
      l_sum_disc_price_dvalid       => PriceSummaryWriter_inst_l_sum_disc_price_dvalid,
      l_sum_disc_price_last         => PriceSummaryWriter_inst_l_sum_disc_price_last,
      l_sum_disc_price              => PriceSummaryWriter_inst_l_sum_disc_price,
      l_sum_charge_valid            => PriceSummaryWriter_inst_l_sum_charge_valid,
      l_sum_charge_ready            => PriceSummaryWriter_inst_l_sum_charge_ready,
      l_sum_charge_dvalid           => PriceSummaryWriter_inst_l_sum_charge_dvalid,
      l_sum_charge_last             => PriceSummaryWriter_inst_l_sum_charge_last,
      l_sum_charge                  => PriceSummaryWriter_inst_l_sum_charge,
      l_avg_qty_valid               => PriceSummaryWriter_inst_l_avg_qty_valid,
      l_avg_qty_ready               => PriceSummaryWriter_inst_l_avg_qty_ready,
      l_avg_qty_dvalid              => PriceSummaryWriter_inst_l_avg_qty_dvalid,
      l_avg_qty_last                => PriceSummaryWriter_inst_l_avg_qty_last,
      l_avg_qty                     => PriceSummaryWriter_inst_l_avg_qty,
      l_avg_price_valid             => PriceSummaryWriter_inst_l_avg_price_valid,
      l_avg_price_ready             => PriceSummaryWriter_inst_l_avg_price_ready,
      l_avg_price_dvalid            => PriceSummaryWriter_inst_l_avg_price_dvalid,
      l_avg_price_last              => PriceSummaryWriter_inst_l_avg_price_last,
      l_avg_price                   => PriceSummaryWriter_inst_l_avg_price,
      l_avg_disc_valid              => PriceSummaryWriter_inst_l_avg_disc_valid,
      l_avg_disc_ready              => PriceSummaryWriter_inst_l_avg_disc_ready,
      l_avg_disc_dvalid             => PriceSummaryWriter_inst_l_avg_disc_dvalid,
      l_avg_disc_last               => PriceSummaryWriter_inst_l_avg_disc_last,
      l_avg_disc                    => PriceSummaryWriter_inst_l_avg_disc,
      l_count_order_valid           => PriceSummaryWriter_inst_l_count_order_valid,
      l_count_order_ready           => PriceSummaryWriter_inst_l_count_order_ready,
      l_count_order_dvalid          => PriceSummaryWriter_inst_l_count_order_dvalid,
      l_count_order_last            => PriceSummaryWriter_inst_l_count_order_last,
      l_count_order                 => PriceSummaryWriter_inst_l_count_order,
      l_returnflag_o_unl_valid      => PriceSummaryWriter_inst_l_returnflag_o_unl_valid,
      l_returnflag_o_unl_ready      => PriceSummaryWriter_inst_l_returnflag_o_unl_ready,
      l_returnflag_o_unl_tag        => PriceSummaryWriter_inst_l_returnflag_o_unl_tag,
      l_linestatus_o_unl_valid      => PriceSummaryWriter_inst_l_linestatus_o_unl_valid,
      l_linestatus_o_unl_ready      => PriceSummaryWriter_inst_l_linestatus_o_unl_ready,
      l_linestatus_o_unl_tag        => PriceSummaryWriter_inst_l_linestatus_o_unl_tag,
      l_sum_qty_unl_valid           => PriceSummaryWriter_inst_l_sum_qty_unl_valid,
      l_sum_qty_unl_ready           => PriceSummaryWriter_inst_l_sum_qty_unl_ready,
      l_sum_qty_unl_tag             => PriceSummaryWriter_inst_l_sum_qty_unl_tag,
      l_sum_base_price_unl_valid    => PriceSummaryWriter_inst_l_sum_base_price_unl_valid,
      l_sum_base_price_unl_ready    => PriceSummaryWriter_inst_l_sum_base_price_unl_ready,
      l_sum_base_price_unl_tag      => PriceSummaryWriter_inst_l_sum_base_price_unl_tag,
      l_sum_disc_price_unl_valid    => PriceSummaryWriter_inst_l_sum_disc_price_unl_valid,
      l_sum_disc_price_unl_ready    => PriceSummaryWriter_inst_l_sum_disc_price_unl_ready,
      l_sum_disc_price_unl_tag      => PriceSummaryWriter_inst_l_sum_disc_price_unl_tag,
      l_sum_charge_unl_valid        => PriceSummaryWriter_inst_l_sum_charge_unl_valid,
      l_sum_charge_unl_ready        => PriceSummaryWriter_inst_l_sum_charge_unl_ready,
      l_sum_charge_unl_tag          => PriceSummaryWriter_inst_l_sum_charge_unl_tag,
      l_avg_qty_unl_valid           => PriceSummaryWriter_inst_l_avg_qty_unl_valid,
      l_avg_qty_unl_ready           => PriceSummaryWriter_inst_l_avg_qty_unl_ready,
      l_avg_qty_unl_tag             => PriceSummaryWriter_inst_l_avg_qty_unl_tag,
      l_avg_price_unl_valid         => PriceSummaryWriter_inst_l_avg_price_unl_valid,
      l_avg_price_unl_ready         => PriceSummaryWriter_inst_l_avg_price_unl_ready,
      l_avg_price_unl_tag           => PriceSummaryWriter_inst_l_avg_price_unl_tag,
      l_avg_disc_unl_valid          => PriceSummaryWriter_inst_l_avg_disc_unl_valid,
      l_avg_disc_unl_ready          => PriceSummaryWriter_inst_l_avg_disc_unl_ready,
      l_avg_disc_unl_tag            => PriceSummaryWriter_inst_l_avg_disc_unl_tag,
      l_count_order_unl_valid       => PriceSummaryWriter_inst_l_count_order_unl_valid,
      l_count_order_unl_ready       => PriceSummaryWriter_inst_l_count_order_unl_ready,
      l_count_order_unl_tag         => PriceSummaryWriter_inst_l_count_order_unl_tag,
      l_returnflag_o_cmd_valid      => PriceSummaryWriter_inst_l_returnflag_o_cmd_valid,
      l_returnflag_o_cmd_ready      => PriceSummaryWriter_inst_l_returnflag_o_cmd_ready,
      l_returnflag_o_cmd_firstIdx   => PriceSummaryWriter_inst_l_returnflag_o_cmd_firstIdx,
      l_returnflag_o_cmd_lastIdx    => PriceSummaryWriter_inst_l_returnflag_o_cmd_lastIdx,
      l_returnflag_o_cmd_tag        => PriceSummaryWriter_inst_l_returnflag_o_cmd_tag,
      l_linestatus_o_cmd_valid      => PriceSummaryWriter_inst_l_linestatus_o_cmd_valid,
      l_linestatus_o_cmd_ready      => PriceSummaryWriter_inst_l_linestatus_o_cmd_ready,
      l_linestatus_o_cmd_firstIdx   => PriceSummaryWriter_inst_l_linestatus_o_cmd_firstIdx,
      l_linestatus_o_cmd_lastIdx    => PriceSummaryWriter_inst_l_linestatus_o_cmd_lastIdx,
      l_linestatus_o_cmd_tag        => PriceSummaryWriter_inst_l_linestatus_o_cmd_tag,
      l_sum_qty_cmd_valid           => PriceSummaryWriter_inst_l_sum_qty_cmd_valid,
      l_sum_qty_cmd_ready           => PriceSummaryWriter_inst_l_sum_qty_cmd_ready,
      l_sum_qty_cmd_firstIdx        => PriceSummaryWriter_inst_l_sum_qty_cmd_firstIdx,
      l_sum_qty_cmd_lastIdx         => PriceSummaryWriter_inst_l_sum_qty_cmd_lastIdx,
      l_sum_qty_cmd_tag             => PriceSummaryWriter_inst_l_sum_qty_cmd_tag,
      l_sum_base_price_cmd_valid    => PriceSummaryWriter_inst_l_sum_base_price_cmd_valid,
      l_sum_base_price_cmd_ready    => PriceSummaryWriter_inst_l_sum_base_price_cmd_ready,
      l_sum_base_price_cmd_firstIdx => PriceSummaryWriter_inst_l_sum_base_price_cmd_firstIdx,
      l_sum_base_price_cmd_lastIdx  => PriceSummaryWriter_inst_l_sum_base_price_cmd_lastIdx,
      l_sum_base_price_cmd_tag      => PriceSummaryWriter_inst_l_sum_base_price_cmd_tag,
      l_sum_disc_price_cmd_valid    => PriceSummaryWriter_inst_l_sum_disc_price_cmd_valid,
      l_sum_disc_price_cmd_ready    => PriceSummaryWriter_inst_l_sum_disc_price_cmd_ready,
      l_sum_disc_price_cmd_firstIdx => PriceSummaryWriter_inst_l_sum_disc_price_cmd_firstIdx,
      l_sum_disc_price_cmd_lastIdx  => PriceSummaryWriter_inst_l_sum_disc_price_cmd_lastIdx,
      l_sum_disc_price_cmd_tag      => PriceSummaryWriter_inst_l_sum_disc_price_cmd_tag,
      l_sum_charge_cmd_valid        => PriceSummaryWriter_inst_l_sum_charge_cmd_valid,
      l_sum_charge_cmd_ready        => PriceSummaryWriter_inst_l_sum_charge_cmd_ready,
      l_sum_charge_cmd_firstIdx     => PriceSummaryWriter_inst_l_sum_charge_cmd_firstIdx,
      l_sum_charge_cmd_lastIdx      => PriceSummaryWriter_inst_l_sum_charge_cmd_lastIdx,
      l_sum_charge_cmd_tag          => PriceSummaryWriter_inst_l_sum_charge_cmd_tag,
      l_avg_qty_cmd_valid           => PriceSummaryWriter_inst_l_avg_qty_cmd_valid,
      l_avg_qty_cmd_ready           => PriceSummaryWriter_inst_l_avg_qty_cmd_ready,
      l_avg_qty_cmd_firstIdx        => PriceSummaryWriter_inst_l_avg_qty_cmd_firstIdx,
      l_avg_qty_cmd_lastIdx         => PriceSummaryWriter_inst_l_avg_qty_cmd_lastIdx,
      l_avg_qty_cmd_tag             => PriceSummaryWriter_inst_l_avg_qty_cmd_tag,
      l_avg_price_cmd_valid         => PriceSummaryWriter_inst_l_avg_price_cmd_valid,
      l_avg_price_cmd_ready         => PriceSummaryWriter_inst_l_avg_price_cmd_ready,
      l_avg_price_cmd_firstIdx      => PriceSummaryWriter_inst_l_avg_price_cmd_firstIdx,
      l_avg_price_cmd_lastIdx       => PriceSummaryWriter_inst_l_avg_price_cmd_lastIdx,
      l_avg_price_cmd_tag           => PriceSummaryWriter_inst_l_avg_price_cmd_tag,
      l_avg_disc_cmd_valid          => PriceSummaryWriter_inst_l_avg_disc_cmd_valid,
      l_avg_disc_cmd_ready          => PriceSummaryWriter_inst_l_avg_disc_cmd_ready,
      l_avg_disc_cmd_firstIdx       => PriceSummaryWriter_inst_l_avg_disc_cmd_firstIdx,
      l_avg_disc_cmd_lastIdx        => PriceSummaryWriter_inst_l_avg_disc_cmd_lastIdx,
      l_avg_disc_cmd_tag            => PriceSummaryWriter_inst_l_avg_disc_cmd_tag,
      l_count_order_cmd_valid       => PriceSummaryWriter_inst_l_count_order_cmd_valid,
      l_count_order_cmd_ready       => PriceSummaryWriter_inst_l_count_order_cmd_ready,
      l_count_order_cmd_firstIdx    => PriceSummaryWriter_inst_l_count_order_cmd_firstIdx,
      l_count_order_cmd_lastIdx     => PriceSummaryWriter_inst_l_count_order_cmd_lastIdx,
      l_count_order_cmd_tag         => PriceSummaryWriter_inst_l_count_order_cmd_tag,
      start                         => PriceSummaryWriter_inst_start,
      stop                          => PriceSummaryWriter_inst_stop,
      reset                         => PriceSummaryWriter_inst_reset,
      idle                          => PriceSummaryWriter_inst_idle,
      busy                          => PriceSummaryWriter_inst_busy,
      done                          => PriceSummaryWriter_inst_done,
      result                        => PriceSummaryWriter_inst_result,
      l_firstidx                    => PriceSummaryWriter_inst_l_firstidx,
      l_lastidx                     => PriceSummaryWriter_inst_l_lastidx
    );

  mmio_inst : mmio
    port map (
      kcd_clk                        => kcd_clk,
      kcd_reset                      => kcd_reset,
      f_start_data                   => mmio_inst_f_start_data,
      f_stop_data                    => mmio_inst_f_stop_data,
      f_reset_data                   => mmio_inst_f_reset_data,
      f_idle_write_data              => mmio_inst_f_idle_write_data,
      f_busy_write_data              => mmio_inst_f_busy_write_data,
      f_done_write_data              => mmio_inst_f_done_write_data,
      f_result_write_data            => mmio_inst_f_result_write_data,
      f_l_firstidx_data              => mmio_inst_f_l_firstidx_data,
      f_l_lastidx_data               => mmio_inst_f_l_lastidx_data,
      f_l_returnflag_o_offsets_data  => mmio_inst_f_l_returnflag_o_offsets_data,
      f_l_returnflag_o_values_data   => mmio_inst_f_l_returnflag_o_values_data,
      f_l_linestatus_o_offsets_data  => mmio_inst_f_l_linestatus_o_offsets_data,
      f_l_linestatus_o_values_data   => mmio_inst_f_l_linestatus_o_values_data,
      f_l_sum_qty_values_data        => mmio_inst_f_l_sum_qty_values_data,
      f_l_sum_base_price_values_data => mmio_inst_f_l_sum_base_price_values_data,
      f_l_sum_disc_price_values_data => mmio_inst_f_l_sum_disc_price_values_data,
      f_l_sum_charge_values_data     => mmio_inst_f_l_sum_charge_values_data,
      f_l_avg_qty_values_data        => mmio_inst_f_l_avg_qty_values_data,
      f_l_avg_price_values_data      => mmio_inst_f_l_avg_price_values_data,
      f_l_avg_disc_values_data       => mmio_inst_f_l_avg_disc_values_data,
      f_l_count_order_values_data    => mmio_inst_f_l_count_order_values_data,
      mmio_awvalid                   => mmio_inst_mmio_awvalid,
      mmio_awready                   => mmio_inst_mmio_awready,
      mmio_awaddr                    => mmio_inst_mmio_awaddr,
      mmio_wvalid                    => mmio_inst_mmio_wvalid,
      mmio_wready                    => mmio_inst_mmio_wready,
      mmio_wdata                     => mmio_inst_mmio_wdata,
      mmio_wstrb                     => mmio_inst_mmio_wstrb,
      mmio_bvalid                    => mmio_inst_mmio_bvalid,
      mmio_bready                    => mmio_inst_mmio_bready,
      mmio_bresp                     => mmio_inst_mmio_bresp,
      mmio_arvalid                   => mmio_inst_mmio_arvalid,
      mmio_arready                   => mmio_inst_mmio_arready,
      mmio_araddr                    => mmio_inst_mmio_araddr,
      mmio_rvalid                    => mmio_inst_mmio_rvalid,
      mmio_rready                    => mmio_inst_mmio_rready,
      mmio_rdata                     => mmio_inst_mmio_rdata,
      mmio_rresp                     => mmio_inst_mmio_rresp
    );

  l_returnflag_o_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 2,
      BUS_ADDR_WIDTH => L_RETURNFLAG_O_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => l_returnflag_o_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => l_returnflag_o_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => l_returnflag_o_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => l_returnflag_o_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => l_returnflag_o_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => l_returnflag_o_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => l_returnflag_o_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => l_returnflag_o_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => l_returnflag_o_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => l_returnflag_o_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => l_returnflag_o_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => l_returnflag_o_cmd_accm_inst_ctrl
    );

  l_linestatus_o_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 2,
      BUS_ADDR_WIDTH => L_LINESTATUS_O_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => l_linestatus_o_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => l_linestatus_o_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => l_linestatus_o_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => l_linestatus_o_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => l_linestatus_o_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => l_linestatus_o_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => l_linestatus_o_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => l_linestatus_o_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => l_linestatus_o_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => l_linestatus_o_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => l_linestatus_o_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => l_linestatus_o_cmd_accm_inst_ctrl
    );

  l_sum_qty_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => L_SUM_QTY_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => l_sum_qty_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => l_sum_qty_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => l_sum_qty_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => l_sum_qty_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => l_sum_qty_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => l_sum_qty_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => l_sum_qty_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => l_sum_qty_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => l_sum_qty_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => l_sum_qty_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => l_sum_qty_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => l_sum_qty_cmd_accm_inst_ctrl
    );

  l_sum_base_price_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => L_SUM_BASE_PRICE_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => l_sum_base_price_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => l_sum_base_price_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => l_sum_base_price_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => l_sum_base_price_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => l_sum_base_price_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => l_sum_base_price_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => l_sum_base_price_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => l_sum_base_price_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => l_sum_base_price_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => l_sum_base_price_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => l_sum_base_price_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => l_sum_base_price_cmd_accm_inst_ctrl
    );

  l_sum_disc_price_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => L_SUM_DISC_PRICE_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => l_sum_disc_price_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => l_sum_disc_price_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => l_sum_disc_price_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => l_sum_disc_price_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => l_sum_disc_price_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => l_sum_disc_price_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => l_sum_disc_price_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => l_sum_disc_price_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => l_sum_disc_price_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => l_sum_disc_price_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => l_sum_disc_price_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => l_sum_disc_price_cmd_accm_inst_ctrl
    );

  l_sum_charge_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => L_SUM_CHARGE_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => l_sum_charge_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => l_sum_charge_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => l_sum_charge_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => l_sum_charge_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => l_sum_charge_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => l_sum_charge_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => l_sum_charge_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => l_sum_charge_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => l_sum_charge_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => l_sum_charge_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => l_sum_charge_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => l_sum_charge_cmd_accm_inst_ctrl
    );

  l_avg_qty_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => L_AVG_QTY_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => l_avg_qty_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => l_avg_qty_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => l_avg_qty_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => l_avg_qty_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => l_avg_qty_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => l_avg_qty_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => l_avg_qty_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => l_avg_qty_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => l_avg_qty_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => l_avg_qty_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => l_avg_qty_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => l_avg_qty_cmd_accm_inst_ctrl
    );

  l_avg_price_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => L_AVG_PRICE_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => l_avg_price_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => l_avg_price_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => l_avg_price_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => l_avg_price_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => l_avg_price_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => l_avg_price_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => l_avg_price_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => l_avg_price_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => l_avg_price_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => l_avg_price_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => l_avg_price_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => l_avg_price_cmd_accm_inst_ctrl
    );

  l_avg_disc_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => L_AVG_DISC_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => l_avg_disc_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => l_avg_disc_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => l_avg_disc_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => l_avg_disc_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => l_avg_disc_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => l_avg_disc_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => l_avg_disc_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => l_avg_disc_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => l_avg_disc_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => l_avg_disc_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => l_avg_disc_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => l_avg_disc_cmd_accm_inst_ctrl
    );

  l_count_order_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => L_COUNT_ORDER_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => l_count_order_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => l_count_order_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => l_count_order_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => l_count_order_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => l_count_order_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => l_count_order_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => l_count_order_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => l_count_order_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => l_count_order_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => l_count_order_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => l_count_order_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => l_count_order_cmd_accm_inst_ctrl
    );

  l_returnflag_o_valid                               <= PriceSummaryWriter_inst_l_returnflag_o_valid;
  PriceSummaryWriter_inst_l_returnflag_o_ready       <= l_returnflag_o_ready;
  l_returnflag_o_dvalid                              <= PriceSummaryWriter_inst_l_returnflag_o_dvalid;
  l_returnflag_o_last                                <= PriceSummaryWriter_inst_l_returnflag_o_last;
  l_returnflag_o_length                              <= PriceSummaryWriter_inst_l_returnflag_o_length;
  l_returnflag_o_count                               <= PriceSummaryWriter_inst_l_returnflag_o_count;
  l_returnflag_o_chars_valid                         <= PriceSummaryWriter_inst_l_returnflag_o_chars_valid;
  PriceSummaryWriter_inst_l_returnflag_o_chars_ready <= l_returnflag_o_chars_ready;
  l_returnflag_o_chars_dvalid                        <= PriceSummaryWriter_inst_l_returnflag_o_chars_dvalid;
  l_returnflag_o_chars_last                          <= PriceSummaryWriter_inst_l_returnflag_o_chars_last;
  l_returnflag_o_chars                               <= PriceSummaryWriter_inst_l_returnflag_o_chars;
  l_returnflag_o_chars_count                         <= PriceSummaryWriter_inst_l_returnflag_o_chars_count;

  l_linestatus_o_valid                               <= PriceSummaryWriter_inst_l_linestatus_o_valid;
  PriceSummaryWriter_inst_l_linestatus_o_ready       <= l_linestatus_o_ready;
  l_linestatus_o_dvalid                              <= PriceSummaryWriter_inst_l_linestatus_o_dvalid;
  l_linestatus_o_last                                <= PriceSummaryWriter_inst_l_linestatus_o_last;
  l_linestatus_o_length                              <= PriceSummaryWriter_inst_l_linestatus_o_length;
  l_linestatus_o_count                               <= PriceSummaryWriter_inst_l_linestatus_o_count;
  l_linestatus_o_chars_valid                         <= PriceSummaryWriter_inst_l_linestatus_o_chars_valid;
  PriceSummaryWriter_inst_l_linestatus_o_chars_ready <= l_linestatus_o_chars_ready;
  l_linestatus_o_chars_dvalid                        <= PriceSummaryWriter_inst_l_linestatus_o_chars_dvalid;
  l_linestatus_o_chars_last                          <= PriceSummaryWriter_inst_l_linestatus_o_chars_last;
  l_linestatus_o_chars                               <= PriceSummaryWriter_inst_l_linestatus_o_chars;
  l_linestatus_o_chars_count                         <= PriceSummaryWriter_inst_l_linestatus_o_chars_count;

  l_sum_qty_valid                                    <= PriceSummaryWriter_inst_l_sum_qty_valid;
  PriceSummaryWriter_inst_l_sum_qty_ready            <= l_sum_qty_ready;
  l_sum_qty_dvalid                                   <= PriceSummaryWriter_inst_l_sum_qty_dvalid;
  l_sum_qty_last                                     <= PriceSummaryWriter_inst_l_sum_qty_last;
  l_sum_qty                                          <= PriceSummaryWriter_inst_l_sum_qty;

  l_sum_base_price_valid                             <= PriceSummaryWriter_inst_l_sum_base_price_valid;
  PriceSummaryWriter_inst_l_sum_base_price_ready     <= l_sum_base_price_ready;
  l_sum_base_price_dvalid                            <= PriceSummaryWriter_inst_l_sum_base_price_dvalid;
  l_sum_base_price_last                              <= PriceSummaryWriter_inst_l_sum_base_price_last;
  l_sum_base_price                                   <= PriceSummaryWriter_inst_l_sum_base_price;

  l_sum_disc_price_valid                             <= PriceSummaryWriter_inst_l_sum_disc_price_valid;
  PriceSummaryWriter_inst_l_sum_disc_price_ready     <= l_sum_disc_price_ready;
  l_sum_disc_price_dvalid                            <= PriceSummaryWriter_inst_l_sum_disc_price_dvalid;
  l_sum_disc_price_last                              <= PriceSummaryWriter_inst_l_sum_disc_price_last;
  l_sum_disc_price                                   <= PriceSummaryWriter_inst_l_sum_disc_price;

  l_sum_charge_valid                                 <= PriceSummaryWriter_inst_l_sum_charge_valid;
  PriceSummaryWriter_inst_l_sum_charge_ready         <= l_sum_charge_ready;
  l_sum_charge_dvalid                                <= PriceSummaryWriter_inst_l_sum_charge_dvalid;
  l_sum_charge_last                                  <= PriceSummaryWriter_inst_l_sum_charge_last;
  l_sum_charge                                       <= PriceSummaryWriter_inst_l_sum_charge;

  l_avg_qty_valid                                    <= PriceSummaryWriter_inst_l_avg_qty_valid;
  PriceSummaryWriter_inst_l_avg_qty_ready            <= l_avg_qty_ready;
  l_avg_qty_dvalid                                   <= PriceSummaryWriter_inst_l_avg_qty_dvalid;
  l_avg_qty_last                                     <= PriceSummaryWriter_inst_l_avg_qty_last;
  l_avg_qty                                          <= PriceSummaryWriter_inst_l_avg_qty;

  l_avg_price_valid                                  <= PriceSummaryWriter_inst_l_avg_price_valid;
  PriceSummaryWriter_inst_l_avg_price_ready          <= l_avg_price_ready;
  l_avg_price_dvalid                                 <= PriceSummaryWriter_inst_l_avg_price_dvalid;
  l_avg_price_last                                   <= PriceSummaryWriter_inst_l_avg_price_last;
  l_avg_price                                        <= PriceSummaryWriter_inst_l_avg_price;

  l_avg_disc_valid                                   <= PriceSummaryWriter_inst_l_avg_disc_valid;
  PriceSummaryWriter_inst_l_avg_disc_ready           <= l_avg_disc_ready;
  l_avg_disc_dvalid                                  <= PriceSummaryWriter_inst_l_avg_disc_dvalid;
  l_avg_disc_last                                    <= PriceSummaryWriter_inst_l_avg_disc_last;
  l_avg_disc                                         <= PriceSummaryWriter_inst_l_avg_disc;

  l_count_order_valid                                <= PriceSummaryWriter_inst_l_count_order_valid;
  PriceSummaryWriter_inst_l_count_order_ready        <= l_count_order_ready;
  l_count_order_dvalid                               <= PriceSummaryWriter_inst_l_count_order_dvalid;
  l_count_order_last                                 <= PriceSummaryWriter_inst_l_count_order_last;
  l_count_order                                      <= PriceSummaryWriter_inst_l_count_order;

  l_returnflag_o_cmd_valid                           <= l_returnflag_o_cmd_accm_inst_nucleus_cmd_valid;
  l_returnflag_o_cmd_accm_inst_nucleus_cmd_ready     <= l_returnflag_o_cmd_ready;
  l_returnflag_o_cmd_firstIdx                        <= l_returnflag_o_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_returnflag_o_cmd_lastIdx                         <= l_returnflag_o_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_returnflag_o_cmd_ctrl                            <= l_returnflag_o_cmd_accm_inst_nucleus_cmd_ctrl;
  l_returnflag_o_cmd_tag                             <= l_returnflag_o_cmd_accm_inst_nucleus_cmd_tag;

  l_linestatus_o_cmd_valid                           <= l_linestatus_o_cmd_accm_inst_nucleus_cmd_valid;
  l_linestatus_o_cmd_accm_inst_nucleus_cmd_ready     <= l_linestatus_o_cmd_ready;
  l_linestatus_o_cmd_firstIdx                        <= l_linestatus_o_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_linestatus_o_cmd_lastIdx                         <= l_linestatus_o_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_linestatus_o_cmd_ctrl                            <= l_linestatus_o_cmd_accm_inst_nucleus_cmd_ctrl;
  l_linestatus_o_cmd_tag                             <= l_linestatus_o_cmd_accm_inst_nucleus_cmd_tag;

  l_sum_qty_cmd_valid                                <= l_sum_qty_cmd_accm_inst_nucleus_cmd_valid;
  l_sum_qty_cmd_accm_inst_nucleus_cmd_ready          <= l_sum_qty_cmd_ready;
  l_sum_qty_cmd_firstIdx                             <= l_sum_qty_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_sum_qty_cmd_lastIdx                              <= l_sum_qty_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_sum_qty_cmd_ctrl                                 <= l_sum_qty_cmd_accm_inst_nucleus_cmd_ctrl;
  l_sum_qty_cmd_tag                                  <= l_sum_qty_cmd_accm_inst_nucleus_cmd_tag;

  l_sum_base_price_cmd_valid                         <= l_sum_base_price_cmd_accm_inst_nucleus_cmd_valid;
  l_sum_base_price_cmd_accm_inst_nucleus_cmd_ready   <= l_sum_base_price_cmd_ready;
  l_sum_base_price_cmd_firstIdx                      <= l_sum_base_price_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_sum_base_price_cmd_lastIdx                       <= l_sum_base_price_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_sum_base_price_cmd_ctrl                          <= l_sum_base_price_cmd_accm_inst_nucleus_cmd_ctrl;
  l_sum_base_price_cmd_tag                           <= l_sum_base_price_cmd_accm_inst_nucleus_cmd_tag;

  l_sum_disc_price_cmd_valid                         <= l_sum_disc_price_cmd_accm_inst_nucleus_cmd_valid;
  l_sum_disc_price_cmd_accm_inst_nucleus_cmd_ready   <= l_sum_disc_price_cmd_ready;
  l_sum_disc_price_cmd_firstIdx                      <= l_sum_disc_price_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_sum_disc_price_cmd_lastIdx                       <= l_sum_disc_price_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_sum_disc_price_cmd_ctrl                          <= l_sum_disc_price_cmd_accm_inst_nucleus_cmd_ctrl;
  l_sum_disc_price_cmd_tag                           <= l_sum_disc_price_cmd_accm_inst_nucleus_cmd_tag;

  l_sum_charge_cmd_valid                             <= l_sum_charge_cmd_accm_inst_nucleus_cmd_valid;
  l_sum_charge_cmd_accm_inst_nucleus_cmd_ready       <= l_sum_charge_cmd_ready;
  l_sum_charge_cmd_firstIdx                          <= l_sum_charge_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_sum_charge_cmd_lastIdx                           <= l_sum_charge_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_sum_charge_cmd_ctrl                              <= l_sum_charge_cmd_accm_inst_nucleus_cmd_ctrl;
  l_sum_charge_cmd_tag                               <= l_sum_charge_cmd_accm_inst_nucleus_cmd_tag;

  l_avg_qty_cmd_valid                                <= l_avg_qty_cmd_accm_inst_nucleus_cmd_valid;
  l_avg_qty_cmd_accm_inst_nucleus_cmd_ready          <= l_avg_qty_cmd_ready;
  l_avg_qty_cmd_firstIdx                             <= l_avg_qty_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_avg_qty_cmd_lastIdx                              <= l_avg_qty_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_avg_qty_cmd_ctrl                                 <= l_avg_qty_cmd_accm_inst_nucleus_cmd_ctrl;
  l_avg_qty_cmd_tag                                  <= l_avg_qty_cmd_accm_inst_nucleus_cmd_tag;

  l_avg_price_cmd_valid                              <= l_avg_price_cmd_accm_inst_nucleus_cmd_valid;
  l_avg_price_cmd_accm_inst_nucleus_cmd_ready        <= l_avg_price_cmd_ready;
  l_avg_price_cmd_firstIdx                           <= l_avg_price_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_avg_price_cmd_lastIdx                            <= l_avg_price_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_avg_price_cmd_ctrl                               <= l_avg_price_cmd_accm_inst_nucleus_cmd_ctrl;
  l_avg_price_cmd_tag                                <= l_avg_price_cmd_accm_inst_nucleus_cmd_tag;

  l_avg_disc_cmd_valid                               <= l_avg_disc_cmd_accm_inst_nucleus_cmd_valid;
  l_avg_disc_cmd_accm_inst_nucleus_cmd_ready         <= l_avg_disc_cmd_ready;
  l_avg_disc_cmd_firstIdx                            <= l_avg_disc_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_avg_disc_cmd_lastIdx                             <= l_avg_disc_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_avg_disc_cmd_ctrl                                <= l_avg_disc_cmd_accm_inst_nucleus_cmd_ctrl;
  l_avg_disc_cmd_tag                                 <= l_avg_disc_cmd_accm_inst_nucleus_cmd_tag;

  l_count_order_cmd_valid                            <= l_count_order_cmd_accm_inst_nucleus_cmd_valid;
  l_count_order_cmd_accm_inst_nucleus_cmd_ready      <= l_count_order_cmd_ready;
  l_count_order_cmd_firstIdx                         <= l_count_order_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_count_order_cmd_lastIdx                          <= l_count_order_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_count_order_cmd_ctrl                             <= l_count_order_cmd_accm_inst_nucleus_cmd_ctrl;
  l_count_order_cmd_tag                              <= l_count_order_cmd_accm_inst_nucleus_cmd_tag;

  PriceSummaryWriter_inst_l_returnflag_o_unl_valid   <= l_returnflag_o_unl_valid;
  l_returnflag_o_unl_ready                           <= PriceSummaryWriter_inst_l_returnflag_o_unl_ready;
  PriceSummaryWriter_inst_l_returnflag_o_unl_tag     <= l_returnflag_o_unl_tag;

  PriceSummaryWriter_inst_l_linestatus_o_unl_valid   <= l_linestatus_o_unl_valid;
  l_linestatus_o_unl_ready                           <= PriceSummaryWriter_inst_l_linestatus_o_unl_ready;
  PriceSummaryWriter_inst_l_linestatus_o_unl_tag     <= l_linestatus_o_unl_tag;

  PriceSummaryWriter_inst_l_sum_qty_unl_valid        <= l_sum_qty_unl_valid;
  l_sum_qty_unl_ready                                <= PriceSummaryWriter_inst_l_sum_qty_unl_ready;
  PriceSummaryWriter_inst_l_sum_qty_unl_tag          <= l_sum_qty_unl_tag;

  PriceSummaryWriter_inst_l_sum_base_price_unl_valid <= l_sum_base_price_unl_valid;
  l_sum_base_price_unl_ready                         <= PriceSummaryWriter_inst_l_sum_base_price_unl_ready;
  PriceSummaryWriter_inst_l_sum_base_price_unl_tag   <= l_sum_base_price_unl_tag;

  PriceSummaryWriter_inst_l_sum_disc_price_unl_valid <= l_sum_disc_price_unl_valid;
  l_sum_disc_price_unl_ready                         <= PriceSummaryWriter_inst_l_sum_disc_price_unl_ready;
  PriceSummaryWriter_inst_l_sum_disc_price_unl_tag   <= l_sum_disc_price_unl_tag;

  PriceSummaryWriter_inst_l_sum_charge_unl_valid     <= l_sum_charge_unl_valid;
  l_sum_charge_unl_ready                             <= PriceSummaryWriter_inst_l_sum_charge_unl_ready;
  PriceSummaryWriter_inst_l_sum_charge_unl_tag       <= l_sum_charge_unl_tag;

  PriceSummaryWriter_inst_l_avg_qty_unl_valid        <= l_avg_qty_unl_valid;
  l_avg_qty_unl_ready                                <= PriceSummaryWriter_inst_l_avg_qty_unl_ready;
  PriceSummaryWriter_inst_l_avg_qty_unl_tag          <= l_avg_qty_unl_tag;

  PriceSummaryWriter_inst_l_avg_price_unl_valid      <= l_avg_price_unl_valid;
  l_avg_price_unl_ready                              <= PriceSummaryWriter_inst_l_avg_price_unl_ready;
  PriceSummaryWriter_inst_l_avg_price_unl_tag        <= l_avg_price_unl_tag;

  PriceSummaryWriter_inst_l_avg_disc_unl_valid       <= l_avg_disc_unl_valid;
  l_avg_disc_unl_ready                               <= PriceSummaryWriter_inst_l_avg_disc_unl_ready;
  PriceSummaryWriter_inst_l_avg_disc_unl_tag         <= l_avg_disc_unl_tag;

  PriceSummaryWriter_inst_l_count_order_unl_valid    <= l_count_order_unl_valid;
  l_count_order_unl_ready                            <= PriceSummaryWriter_inst_l_count_order_unl_ready;
  PriceSummaryWriter_inst_l_count_order_unl_tag      <= l_count_order_unl_tag;

  PriceSummaryWriter_inst_start                      <= mmio_inst_f_start_data;
  PriceSummaryWriter_inst_stop                       <= mmio_inst_f_stop_data;
  PriceSummaryWriter_inst_reset                      <= mmio_inst_f_reset_data;
  PriceSummaryWriter_inst_l_firstidx                 <= mmio_inst_f_l_firstidx_data;
  PriceSummaryWriter_inst_l_lastidx                  <= mmio_inst_f_l_lastidx_data;
  mmio_inst_f_idle_write_data                        <= PriceSummaryWriter_inst_idle;
  mmio_inst_f_busy_write_data                        <= PriceSummaryWriter_inst_busy;
  mmio_inst_f_done_write_data                        <= PriceSummaryWriter_inst_done;
  mmio_inst_f_result_write_data                      <= PriceSummaryWriter_inst_result;
  mmio_inst_mmio_awvalid                             <= mmio_awvalid;
  mmio_awready                                       <= mmio_inst_mmio_awready;
  mmio_inst_mmio_awaddr                              <= mmio_awaddr;
  mmio_inst_mmio_wvalid                              <= mmio_wvalid;
  mmio_wready                                        <= mmio_inst_mmio_wready;
  mmio_inst_mmio_wdata                               <= mmio_wdata;
  mmio_inst_mmio_wstrb                               <= mmio_wstrb;
  mmio_bvalid                                        <= mmio_inst_mmio_bvalid;
  mmio_inst_mmio_bready                              <= mmio_bready;
  mmio_bresp                                         <= mmio_inst_mmio_bresp;
  mmio_inst_mmio_arvalid                             <= mmio_arvalid;
  mmio_arready                                       <= mmio_inst_mmio_arready;
  mmio_inst_mmio_araddr                              <= mmio_araddr;
  mmio_rvalid                                        <= mmio_inst_mmio_rvalid;
  mmio_inst_mmio_rready                              <= mmio_rready;
  mmio_rdata                                         <= mmio_inst_mmio_rdata;
  mmio_rresp                                         <= mmio_inst_mmio_rresp;

  l_returnflag_o_cmd_accm_inst_kernel_cmd_valid      <= PriceSummaryWriter_inst_l_returnflag_o_cmd_valid;
  PriceSummaryWriter_inst_l_returnflag_o_cmd_ready   <= l_returnflag_o_cmd_accm_inst_kernel_cmd_ready;
  l_returnflag_o_cmd_accm_inst_kernel_cmd_firstIdx   <= PriceSummaryWriter_inst_l_returnflag_o_cmd_firstIdx;
  l_returnflag_o_cmd_accm_inst_kernel_cmd_lastIdx    <= PriceSummaryWriter_inst_l_returnflag_o_cmd_lastIdx;
  l_returnflag_o_cmd_accm_inst_kernel_cmd_tag        <= PriceSummaryWriter_inst_l_returnflag_o_cmd_tag;

  l_linestatus_o_cmd_accm_inst_kernel_cmd_valid      <= PriceSummaryWriter_inst_l_linestatus_o_cmd_valid;
  PriceSummaryWriter_inst_l_linestatus_o_cmd_ready   <= l_linestatus_o_cmd_accm_inst_kernel_cmd_ready;
  l_linestatus_o_cmd_accm_inst_kernel_cmd_firstIdx   <= PriceSummaryWriter_inst_l_linestatus_o_cmd_firstIdx;
  l_linestatus_o_cmd_accm_inst_kernel_cmd_lastIdx    <= PriceSummaryWriter_inst_l_linestatus_o_cmd_lastIdx;
  l_linestatus_o_cmd_accm_inst_kernel_cmd_tag        <= PriceSummaryWriter_inst_l_linestatus_o_cmd_tag;

  l_sum_qty_cmd_accm_inst_kernel_cmd_valid           <= PriceSummaryWriter_inst_l_sum_qty_cmd_valid;
  PriceSummaryWriter_inst_l_sum_qty_cmd_ready        <= l_sum_qty_cmd_accm_inst_kernel_cmd_ready;
  l_sum_qty_cmd_accm_inst_kernel_cmd_firstIdx        <= PriceSummaryWriter_inst_l_sum_qty_cmd_firstIdx;
  l_sum_qty_cmd_accm_inst_kernel_cmd_lastIdx         <= PriceSummaryWriter_inst_l_sum_qty_cmd_lastIdx;
  l_sum_qty_cmd_accm_inst_kernel_cmd_tag             <= PriceSummaryWriter_inst_l_sum_qty_cmd_tag;

  l_sum_base_price_cmd_accm_inst_kernel_cmd_valid    <= PriceSummaryWriter_inst_l_sum_base_price_cmd_valid;
  PriceSummaryWriter_inst_l_sum_base_price_cmd_ready <= l_sum_base_price_cmd_accm_inst_kernel_cmd_ready;
  l_sum_base_price_cmd_accm_inst_kernel_cmd_firstIdx <= PriceSummaryWriter_inst_l_sum_base_price_cmd_firstIdx;
  l_sum_base_price_cmd_accm_inst_kernel_cmd_lastIdx  <= PriceSummaryWriter_inst_l_sum_base_price_cmd_lastIdx;
  l_sum_base_price_cmd_accm_inst_kernel_cmd_tag      <= PriceSummaryWriter_inst_l_sum_base_price_cmd_tag;

  l_sum_disc_price_cmd_accm_inst_kernel_cmd_valid    <= PriceSummaryWriter_inst_l_sum_disc_price_cmd_valid;
  PriceSummaryWriter_inst_l_sum_disc_price_cmd_ready <= l_sum_disc_price_cmd_accm_inst_kernel_cmd_ready;
  l_sum_disc_price_cmd_accm_inst_kernel_cmd_firstIdx <= PriceSummaryWriter_inst_l_sum_disc_price_cmd_firstIdx;
  l_sum_disc_price_cmd_accm_inst_kernel_cmd_lastIdx  <= PriceSummaryWriter_inst_l_sum_disc_price_cmd_lastIdx;
  l_sum_disc_price_cmd_accm_inst_kernel_cmd_tag      <= PriceSummaryWriter_inst_l_sum_disc_price_cmd_tag;

  l_sum_charge_cmd_accm_inst_kernel_cmd_valid        <= PriceSummaryWriter_inst_l_sum_charge_cmd_valid;
  PriceSummaryWriter_inst_l_sum_charge_cmd_ready     <= l_sum_charge_cmd_accm_inst_kernel_cmd_ready;
  l_sum_charge_cmd_accm_inst_kernel_cmd_firstIdx     <= PriceSummaryWriter_inst_l_sum_charge_cmd_firstIdx;
  l_sum_charge_cmd_accm_inst_kernel_cmd_lastIdx      <= PriceSummaryWriter_inst_l_sum_charge_cmd_lastIdx;
  l_sum_charge_cmd_accm_inst_kernel_cmd_tag          <= PriceSummaryWriter_inst_l_sum_charge_cmd_tag;

  l_avg_qty_cmd_accm_inst_kernel_cmd_valid           <= PriceSummaryWriter_inst_l_avg_qty_cmd_valid;
  PriceSummaryWriter_inst_l_avg_qty_cmd_ready        <= l_avg_qty_cmd_accm_inst_kernel_cmd_ready;
  l_avg_qty_cmd_accm_inst_kernel_cmd_firstIdx        <= PriceSummaryWriter_inst_l_avg_qty_cmd_firstIdx;
  l_avg_qty_cmd_accm_inst_kernel_cmd_lastIdx         <= PriceSummaryWriter_inst_l_avg_qty_cmd_lastIdx;
  l_avg_qty_cmd_accm_inst_kernel_cmd_tag             <= PriceSummaryWriter_inst_l_avg_qty_cmd_tag;

  l_avg_price_cmd_accm_inst_kernel_cmd_valid         <= PriceSummaryWriter_inst_l_avg_price_cmd_valid;
  PriceSummaryWriter_inst_l_avg_price_cmd_ready      <= l_avg_price_cmd_accm_inst_kernel_cmd_ready;
  l_avg_price_cmd_accm_inst_kernel_cmd_firstIdx      <= PriceSummaryWriter_inst_l_avg_price_cmd_firstIdx;
  l_avg_price_cmd_accm_inst_kernel_cmd_lastIdx       <= PriceSummaryWriter_inst_l_avg_price_cmd_lastIdx;
  l_avg_price_cmd_accm_inst_kernel_cmd_tag           <= PriceSummaryWriter_inst_l_avg_price_cmd_tag;

  l_avg_disc_cmd_accm_inst_kernel_cmd_valid          <= PriceSummaryWriter_inst_l_avg_disc_cmd_valid;
  PriceSummaryWriter_inst_l_avg_disc_cmd_ready       <= l_avg_disc_cmd_accm_inst_kernel_cmd_ready;
  l_avg_disc_cmd_accm_inst_kernel_cmd_firstIdx       <= PriceSummaryWriter_inst_l_avg_disc_cmd_firstIdx;
  l_avg_disc_cmd_accm_inst_kernel_cmd_lastIdx        <= PriceSummaryWriter_inst_l_avg_disc_cmd_lastIdx;
  l_avg_disc_cmd_accm_inst_kernel_cmd_tag            <= PriceSummaryWriter_inst_l_avg_disc_cmd_tag;

  l_count_order_cmd_accm_inst_kernel_cmd_valid       <= PriceSummaryWriter_inst_l_count_order_cmd_valid;
  PriceSummaryWriter_inst_l_count_order_cmd_ready    <= l_count_order_cmd_accm_inst_kernel_cmd_ready;
  l_count_order_cmd_accm_inst_kernel_cmd_firstIdx    <= PriceSummaryWriter_inst_l_count_order_cmd_firstIdx;
  l_count_order_cmd_accm_inst_kernel_cmd_lastIdx     <= PriceSummaryWriter_inst_l_count_order_cmd_lastIdx;
  l_count_order_cmd_accm_inst_kernel_cmd_tag         <= PriceSummaryWriter_inst_l_count_order_cmd_tag;

  l_returnflag_o_cmd_accm_inst_ctrl(63 downto 0)   <= mmio_inst_f_l_returnflag_o_offsets_data;
  l_returnflag_o_cmd_accm_inst_ctrl(127 downto 64) <= mmio_inst_f_l_returnflag_o_values_data;

  l_linestatus_o_cmd_accm_inst_ctrl(63 downto 0)   <= mmio_inst_f_l_linestatus_o_offsets_data;
  l_linestatus_o_cmd_accm_inst_ctrl(127 downto 64) <= mmio_inst_f_l_linestatus_o_values_data;

  l_sum_qty_cmd_accm_inst_ctrl(63 downto 0)        <= mmio_inst_f_l_sum_qty_values_data;
  l_sum_base_price_cmd_accm_inst_ctrl(63 downto 0) <= mmio_inst_f_l_sum_base_price_values_data;
  l_sum_disc_price_cmd_accm_inst_ctrl(63 downto 0) <= mmio_inst_f_l_sum_disc_price_values_data;
  l_sum_charge_cmd_accm_inst_ctrl(63 downto 0)     <= mmio_inst_f_l_sum_charge_values_data;
  l_avg_qty_cmd_accm_inst_ctrl(63 downto 0)        <= mmio_inst_f_l_avg_qty_values_data;
  l_avg_price_cmd_accm_inst_ctrl(63 downto 0)      <= mmio_inst_f_l_avg_price_values_data;
  l_avg_disc_cmd_accm_inst_ctrl(63 downto 0)       <= mmio_inst_f_l_avg_disc_values_data;
  l_count_order_cmd_accm_inst_ctrl(63 downto 0)    <= mmio_inst_f_l_count_order_values_data;

end architecture;
