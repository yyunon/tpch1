-- Copyright 2018-2019 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
-- This file was generated by Fletchgen. Modify this file at your own risk.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.Interconnect_pkg.all;

entity PriceSummaryWriter_Mantle is
  generic (
    INDEX_WIDTH        : integer := 32;
    TAG_WIDTH          : integer := 1;
    BUS_ADDR_WIDTH     : integer := 64;
    BUS_DATA_WIDTH     : integer := 512;
    BUS_LEN_WIDTH      : integer := 8;
    BUS_BURST_STEP_LEN : integer := 1;
    BUS_BURST_MAX_LEN  : integer := 16
  );
  port (
    bcd_clk            : in  std_logic;
    bcd_reset          : in  std_logic;
    kcd_clk            : in  std_logic;
    kcd_reset          : in  std_logic;
    mmio_awvalid       : in  std_logic;
    mmio_awready       : out std_logic;
    mmio_awaddr        : in  std_logic_vector(31 downto 0);
    mmio_wvalid        : in  std_logic;
    mmio_wready        : out std_logic;
    mmio_wdata         : in  std_logic_vector(31 downto 0);
    mmio_wstrb         : in  std_logic_vector(3 downto 0);
    mmio_bvalid        : out std_logic;
    mmio_bready        : in  std_logic;
    mmio_bresp         : out std_logic_vector(1 downto 0);
    mmio_arvalid       : in  std_logic;
    mmio_arready       : out std_logic;
    mmio_araddr        : in  std_logic_vector(31 downto 0);
    mmio_rvalid        : out std_logic;
    mmio_rready        : in  std_logic;
    mmio_rdata         : out std_logic_vector(31 downto 0);
    mmio_rresp         : out std_logic_vector(1 downto 0);
    wr_mst_wreq_valid  : out std_logic;
    wr_mst_wreq_ready  : in  std_logic;
    wr_mst_wreq_addr   : out std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
    wr_mst_wreq_len    : out std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
    wr_mst_wdat_valid  : out std_logic;
    wr_mst_wdat_ready  : in  std_logic;
    wr_mst_wdat_data   : out std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
    wr_mst_wdat_strobe : out std_logic_vector(BUS_DATA_WIDTH/8-1 downto 0);
    wr_mst_wdat_last   : out std_logic
  );
end entity;

architecture Implementation of PriceSummaryWriter_Mantle is
  component PriceSummaryWriter_Nucleus is
    generic (
      INDEX_WIDTH                     : integer := 32;
      TAG_WIDTH                       : integer := 1;
      L_RETURNFLAG_O_BUS_ADDR_WIDTH   : integer := 64;
      L_LINESTATUS_O_BUS_ADDR_WIDTH   : integer := 64;
      L_SUM_QTY_BUS_ADDR_WIDTH        : integer := 64;
      L_SUM_BASE_PRICE_BUS_ADDR_WIDTH : integer := 64;
      L_SUM_DISC_PRICE_BUS_ADDR_WIDTH : integer := 64;
      L_SUM_CHARGE_BUS_ADDR_WIDTH     : integer := 64;
      L_AVG_QTY_BUS_ADDR_WIDTH        : integer := 64;
      L_AVG_PRICE_BUS_ADDR_WIDTH      : integer := 64;
      L_AVG_DISC_BUS_ADDR_WIDTH       : integer := 64;
      L_COUNT_ORDER_BUS_ADDR_WIDTH    : integer := 64
    );
    port (
      kcd_clk                       : in  std_logic;
      kcd_reset                     : in  std_logic;
      mmio_awvalid                  : in  std_logic;
      mmio_awready                  : out std_logic;
      mmio_awaddr                   : in  std_logic_vector(31 downto 0);
      mmio_wvalid                   : in  std_logic;
      mmio_wready                   : out std_logic;
      mmio_wdata                    : in  std_logic_vector(31 downto 0);
      mmio_wstrb                    : in  std_logic_vector(3 downto 0);
      mmio_bvalid                   : out std_logic;
      mmio_bready                   : in  std_logic;
      mmio_bresp                    : out std_logic_vector(1 downto 0);
      mmio_arvalid                  : in  std_logic;
      mmio_arready                  : out std_logic;
      mmio_araddr                   : in  std_logic_vector(31 downto 0);
      mmio_rvalid                   : out std_logic;
      mmio_rready                   : in  std_logic;
      mmio_rdata                    : out std_logic_vector(31 downto 0);
      mmio_rresp                    : out std_logic_vector(1 downto 0);
      l_returnflag_o_valid          : out std_logic;
      l_returnflag_o_ready          : in  std_logic;
      l_returnflag_o_dvalid         : out std_logic;
      l_returnflag_o_last           : out std_logic;
      l_returnflag_o_length         : out std_logic_vector(31 downto 0);
      l_returnflag_o_count          : out std_logic_vector(0 downto 0);
      l_returnflag_o_chars_valid    : out std_logic;
      l_returnflag_o_chars_ready    : in  std_logic;
      l_returnflag_o_chars_dvalid   : out std_logic;
      l_returnflag_o_chars_last     : out std_logic;
      l_returnflag_o_chars          : out std_logic_vector(7 downto 0);
      l_returnflag_o_chars_count    : out std_logic_vector(0 downto 0);
      l_linestatus_o_valid          : out std_logic;
      l_linestatus_o_ready          : in  std_logic;
      l_linestatus_o_dvalid         : out std_logic;
      l_linestatus_o_last           : out std_logic;
      l_linestatus_o_length         : out std_logic_vector(31 downto 0);
      l_linestatus_o_count          : out std_logic_vector(0 downto 0);
      l_linestatus_o_chars_valid    : out std_logic;
      l_linestatus_o_chars_ready    : in  std_logic;
      l_linestatus_o_chars_dvalid   : out std_logic;
      l_linestatus_o_chars_last     : out std_logic;
      l_linestatus_o_chars          : out std_logic_vector(7 downto 0);
      l_linestatus_o_chars_count    : out std_logic_vector(0 downto 0);
      l_sum_qty_valid               : out std_logic;
      l_sum_qty_ready               : in  std_logic;
      l_sum_qty_dvalid              : out std_logic;
      l_sum_qty_last                : out std_logic;
      l_sum_qty                     : out std_logic_vector(63 downto 0);
      l_sum_base_price_valid        : out std_logic;
      l_sum_base_price_ready        : in  std_logic;
      l_sum_base_price_dvalid       : out std_logic;
      l_sum_base_price_last         : out std_logic;
      l_sum_base_price              : out std_logic_vector(63 downto 0);
      l_sum_disc_price_valid        : out std_logic;
      l_sum_disc_price_ready        : in  std_logic;
      l_sum_disc_price_dvalid       : out std_logic;
      l_sum_disc_price_last         : out std_logic;
      l_sum_disc_price              : out std_logic_vector(63 downto 0);
      l_sum_charge_valid            : out std_logic;
      l_sum_charge_ready            : in  std_logic;
      l_sum_charge_dvalid           : out std_logic;
      l_sum_charge_last             : out std_logic;
      l_sum_charge                  : out std_logic_vector(63 downto 0);
      l_avg_qty_valid               : out std_logic;
      l_avg_qty_ready               : in  std_logic;
      l_avg_qty_dvalid              : out std_logic;
      l_avg_qty_last                : out std_logic;
      l_avg_qty                     : out std_logic_vector(63 downto 0);
      l_avg_price_valid             : out std_logic;
      l_avg_price_ready             : in  std_logic;
      l_avg_price_dvalid            : out std_logic;
      l_avg_price_last              : out std_logic;
      l_avg_price                   : out std_logic_vector(63 downto 0);
      l_avg_disc_valid              : out std_logic;
      l_avg_disc_ready              : in  std_logic;
      l_avg_disc_dvalid             : out std_logic;
      l_avg_disc_last               : out std_logic;
      l_avg_disc                    : out std_logic_vector(63 downto 0);
      l_count_order_valid           : out std_logic;
      l_count_order_ready           : in  std_logic;
      l_count_order_dvalid          : out std_logic;
      l_count_order_last            : out std_logic;
      l_count_order                 : out std_logic_vector(63 downto 0);
      l_returnflag_o_unl_valid      : in  std_logic;
      l_returnflag_o_unl_ready      : out std_logic;
      l_returnflag_o_unl_tag        : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_linestatus_o_unl_valid      : in  std_logic;
      l_linestatus_o_unl_ready      : out std_logic;
      l_linestatus_o_unl_tag        : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_sum_qty_unl_valid           : in  std_logic;
      l_sum_qty_unl_ready           : out std_logic;
      l_sum_qty_unl_tag             : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_sum_base_price_unl_valid    : in  std_logic;
      l_sum_base_price_unl_ready    : out std_logic;
      l_sum_base_price_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_sum_disc_price_unl_valid    : in  std_logic;
      l_sum_disc_price_unl_ready    : out std_logic;
      l_sum_disc_price_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_sum_charge_unl_valid        : in  std_logic;
      l_sum_charge_unl_ready        : out std_logic;
      l_sum_charge_unl_tag          : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_avg_qty_unl_valid           : in  std_logic;
      l_avg_qty_unl_ready           : out std_logic;
      l_avg_qty_unl_tag             : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_avg_price_unl_valid         : in  std_logic;
      l_avg_price_unl_ready         : out std_logic;
      l_avg_price_unl_tag           : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_avg_disc_unl_valid          : in  std_logic;
      l_avg_disc_unl_ready          : out std_logic;
      l_avg_disc_unl_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_count_order_unl_valid       : in  std_logic;
      l_count_order_unl_ready       : out std_logic;
      l_count_order_unl_tag         : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_returnflag_o_cmd_valid      : out std_logic;
      l_returnflag_o_cmd_ready      : in  std_logic;
      l_returnflag_o_cmd_firstIdx   : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_returnflag_o_cmd_lastIdx    : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_returnflag_o_cmd_ctrl       : out std_logic_vector(L_RETURNFLAG_O_BUS_ADDR_WIDTH*2-1 downto 0);
      l_returnflag_o_cmd_tag        : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_linestatus_o_cmd_valid      : out std_logic;
      l_linestatus_o_cmd_ready      : in  std_logic;
      l_linestatus_o_cmd_firstIdx   : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_linestatus_o_cmd_lastIdx    : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_linestatus_o_cmd_ctrl       : out std_logic_vector(L_LINESTATUS_O_BUS_ADDR_WIDTH*2-1 downto 0);
      l_linestatus_o_cmd_tag        : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_sum_qty_cmd_valid           : out std_logic;
      l_sum_qty_cmd_ready           : in  std_logic;
      l_sum_qty_cmd_firstIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_sum_qty_cmd_lastIdx         : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_sum_qty_cmd_ctrl            : out std_logic_vector(L_SUM_QTY_BUS_ADDR_WIDTH-1 downto 0);
      l_sum_qty_cmd_tag             : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_sum_base_price_cmd_valid    : out std_logic;
      l_sum_base_price_cmd_ready    : in  std_logic;
      l_sum_base_price_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_sum_base_price_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_sum_base_price_cmd_ctrl     : out std_logic_vector(L_SUM_BASE_PRICE_BUS_ADDR_WIDTH-1 downto 0);
      l_sum_base_price_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_sum_disc_price_cmd_valid    : out std_logic;
      l_sum_disc_price_cmd_ready    : in  std_logic;
      l_sum_disc_price_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_sum_disc_price_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_sum_disc_price_cmd_ctrl     : out std_logic_vector(L_SUM_DISC_PRICE_BUS_ADDR_WIDTH-1 downto 0);
      l_sum_disc_price_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_sum_charge_cmd_valid        : out std_logic;
      l_sum_charge_cmd_ready        : in  std_logic;
      l_sum_charge_cmd_firstIdx     : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_sum_charge_cmd_lastIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_sum_charge_cmd_ctrl         : out std_logic_vector(L_SUM_CHARGE_BUS_ADDR_WIDTH-1 downto 0);
      l_sum_charge_cmd_tag          : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_avg_qty_cmd_valid           : out std_logic;
      l_avg_qty_cmd_ready           : in  std_logic;
      l_avg_qty_cmd_firstIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_avg_qty_cmd_lastIdx         : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_avg_qty_cmd_ctrl            : out std_logic_vector(L_AVG_QTY_BUS_ADDR_WIDTH-1 downto 0);
      l_avg_qty_cmd_tag             : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_avg_price_cmd_valid         : out std_logic;
      l_avg_price_cmd_ready         : in  std_logic;
      l_avg_price_cmd_firstIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_avg_price_cmd_lastIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_avg_price_cmd_ctrl          : out std_logic_vector(L_AVG_PRICE_BUS_ADDR_WIDTH-1 downto 0);
      l_avg_price_cmd_tag           : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_avg_disc_cmd_valid          : out std_logic;
      l_avg_disc_cmd_ready          : in  std_logic;
      l_avg_disc_cmd_firstIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_avg_disc_cmd_lastIdx        : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_avg_disc_cmd_ctrl           : out std_logic_vector(L_AVG_DISC_BUS_ADDR_WIDTH-1 downto 0);
      l_avg_disc_cmd_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_count_order_cmd_valid       : out std_logic;
      l_count_order_cmd_ready       : in  std_logic;
      l_count_order_cmd_firstIdx    : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_count_order_cmd_lastIdx     : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_count_order_cmd_ctrl        : out std_logic_vector(L_COUNT_ORDER_BUS_ADDR_WIDTH-1 downto 0);
      l_count_order_cmd_tag         : out std_logic_vector(TAG_WIDTH-1 downto 0)
    );
  end component;

  component PriceSummaryWriter_l is
    generic (
      INDEX_WIDTH                         : integer := 32;
      TAG_WIDTH                           : integer := 1;
      L_RETURNFLAG_O_BUS_ADDR_WIDTH       : integer := 64;
      L_RETURNFLAG_O_BUS_DATA_WIDTH       : integer := 512;
      L_RETURNFLAG_O_BUS_LEN_WIDTH        : integer := 8;
      L_RETURNFLAG_O_BUS_BURST_STEP_LEN   : integer := 1;
      L_RETURNFLAG_O_BUS_BURST_MAX_LEN    : integer := 16;
      L_LINESTATUS_O_BUS_ADDR_WIDTH       : integer := 64;
      L_LINESTATUS_O_BUS_DATA_WIDTH       : integer := 512;
      L_LINESTATUS_O_BUS_LEN_WIDTH        : integer := 8;
      L_LINESTATUS_O_BUS_BURST_STEP_LEN   : integer := 1;
      L_LINESTATUS_O_BUS_BURST_MAX_LEN    : integer := 16;
      L_SUM_QTY_BUS_ADDR_WIDTH            : integer := 64;
      L_SUM_QTY_BUS_DATA_WIDTH            : integer := 512;
      L_SUM_QTY_BUS_LEN_WIDTH             : integer := 8;
      L_SUM_QTY_BUS_BURST_STEP_LEN        : integer := 1;
      L_SUM_QTY_BUS_BURST_MAX_LEN         : integer := 16;
      L_SUM_BASE_PRICE_BUS_ADDR_WIDTH     : integer := 64;
      L_SUM_BASE_PRICE_BUS_DATA_WIDTH     : integer := 512;
      L_SUM_BASE_PRICE_BUS_LEN_WIDTH      : integer := 8;
      L_SUM_BASE_PRICE_BUS_BURST_STEP_LEN : integer := 1;
      L_SUM_BASE_PRICE_BUS_BURST_MAX_LEN  : integer := 16;
      L_SUM_DISC_PRICE_BUS_ADDR_WIDTH     : integer := 64;
      L_SUM_DISC_PRICE_BUS_DATA_WIDTH     : integer := 512;
      L_SUM_DISC_PRICE_BUS_LEN_WIDTH      : integer := 8;
      L_SUM_DISC_PRICE_BUS_BURST_STEP_LEN : integer := 1;
      L_SUM_DISC_PRICE_BUS_BURST_MAX_LEN  : integer := 16;
      L_SUM_CHARGE_BUS_ADDR_WIDTH         : integer := 64;
      L_SUM_CHARGE_BUS_DATA_WIDTH         : integer := 512;
      L_SUM_CHARGE_BUS_LEN_WIDTH          : integer := 8;
      L_SUM_CHARGE_BUS_BURST_STEP_LEN     : integer := 1;
      L_SUM_CHARGE_BUS_BURST_MAX_LEN      : integer := 16;
      L_AVG_QTY_BUS_ADDR_WIDTH            : integer := 64;
      L_AVG_QTY_BUS_DATA_WIDTH            : integer := 512;
      L_AVG_QTY_BUS_LEN_WIDTH             : integer := 8;
      L_AVG_QTY_BUS_BURST_STEP_LEN        : integer := 1;
      L_AVG_QTY_BUS_BURST_MAX_LEN         : integer := 16;
      L_AVG_PRICE_BUS_ADDR_WIDTH          : integer := 64;
      L_AVG_PRICE_BUS_DATA_WIDTH          : integer := 512;
      L_AVG_PRICE_BUS_LEN_WIDTH           : integer := 8;
      L_AVG_PRICE_BUS_BURST_STEP_LEN      : integer := 1;
      L_AVG_PRICE_BUS_BURST_MAX_LEN       : integer := 16;
      L_AVG_DISC_BUS_ADDR_WIDTH           : integer := 64;
      L_AVG_DISC_BUS_DATA_WIDTH           : integer := 512;
      L_AVG_DISC_BUS_LEN_WIDTH            : integer := 8;
      L_AVG_DISC_BUS_BURST_STEP_LEN       : integer := 1;
      L_AVG_DISC_BUS_BURST_MAX_LEN        : integer := 16;
      L_COUNT_ORDER_BUS_ADDR_WIDTH        : integer := 64;
      L_COUNT_ORDER_BUS_DATA_WIDTH        : integer := 512;
      L_COUNT_ORDER_BUS_LEN_WIDTH         : integer := 8;
      L_COUNT_ORDER_BUS_BURST_STEP_LEN    : integer := 1;
      L_COUNT_ORDER_BUS_BURST_MAX_LEN     : integer := 16
    );
    port (
      bcd_clk                          : in  std_logic;
      bcd_reset                        : in  std_logic;
      kcd_clk                          : in  std_logic;
      kcd_reset                        : in  std_logic;
      l_returnflag_o_valid             : in  std_logic;
      l_returnflag_o_ready             : out std_logic;
      l_returnflag_o_dvalid            : in  std_logic;
      l_returnflag_o_last              : in  std_logic;
      l_returnflag_o_length            : in  std_logic_vector(31 downto 0);
      l_returnflag_o_count             : in  std_logic_vector(0 downto 0);
      l_returnflag_o_chars_valid       : in  std_logic;
      l_returnflag_o_chars_ready       : out std_logic;
      l_returnflag_o_chars_dvalid      : in  std_logic;
      l_returnflag_o_chars_last        : in  std_logic;
      l_returnflag_o_chars             : in  std_logic_vector(7 downto 0);
      l_returnflag_o_chars_count       : in  std_logic_vector(0 downto 0);
      l_returnflag_o_bus_wreq_valid    : out std_logic;
      l_returnflag_o_bus_wreq_ready    : in  std_logic;
      l_returnflag_o_bus_wreq_addr     : out std_logic_vector(L_RETURNFLAG_O_BUS_ADDR_WIDTH-1 downto 0);
      l_returnflag_o_bus_wreq_len      : out std_logic_vector(L_RETURNFLAG_O_BUS_LEN_WIDTH-1 downto 0);
      l_returnflag_o_bus_wdat_valid    : out std_logic;
      l_returnflag_o_bus_wdat_ready    : in  std_logic;
      l_returnflag_o_bus_wdat_data     : out std_logic_vector(L_RETURNFLAG_O_BUS_DATA_WIDTH-1 downto 0);
      l_returnflag_o_bus_wdat_strobe   : out std_logic_vector(L_RETURNFLAG_O_BUS_DATA_WIDTH/8-1 downto 0);
      l_returnflag_o_bus_wdat_last     : out std_logic;
      l_returnflag_o_cmd_valid         : in  std_logic;
      l_returnflag_o_cmd_ready         : out std_logic;
      l_returnflag_o_cmd_firstIdx      : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_returnflag_o_cmd_lastIdx       : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_returnflag_o_cmd_ctrl          : in  std_logic_vector(L_RETURNFLAG_O_BUS_ADDR_WIDTH*2-1 downto 0);
      l_returnflag_o_cmd_tag           : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_returnflag_o_unl_valid         : out std_logic;
      l_returnflag_o_unl_ready         : in  std_logic;
      l_returnflag_o_unl_tag           : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_linestatus_o_valid             : in  std_logic;
      l_linestatus_o_ready             : out std_logic;
      l_linestatus_o_dvalid            : in  std_logic;
      l_linestatus_o_last              : in  std_logic;
      l_linestatus_o_length            : in  std_logic_vector(31 downto 0);
      l_linestatus_o_count             : in  std_logic_vector(0 downto 0);
      l_linestatus_o_chars_valid       : in  std_logic;
      l_linestatus_o_chars_ready       : out std_logic;
      l_linestatus_o_chars_dvalid      : in  std_logic;
      l_linestatus_o_chars_last        : in  std_logic;
      l_linestatus_o_chars             : in  std_logic_vector(7 downto 0);
      l_linestatus_o_chars_count       : in  std_logic_vector(0 downto 0);
      l_linestatus_o_bus_wreq_valid    : out std_logic;
      l_linestatus_o_bus_wreq_ready    : in  std_logic;
      l_linestatus_o_bus_wreq_addr     : out std_logic_vector(L_LINESTATUS_O_BUS_ADDR_WIDTH-1 downto 0);
      l_linestatus_o_bus_wreq_len      : out std_logic_vector(L_LINESTATUS_O_BUS_LEN_WIDTH-1 downto 0);
      l_linestatus_o_bus_wdat_valid    : out std_logic;
      l_linestatus_o_bus_wdat_ready    : in  std_logic;
      l_linestatus_o_bus_wdat_data     : out std_logic_vector(L_LINESTATUS_O_BUS_DATA_WIDTH-1 downto 0);
      l_linestatus_o_bus_wdat_strobe   : out std_logic_vector(L_LINESTATUS_O_BUS_DATA_WIDTH/8-1 downto 0);
      l_linestatus_o_bus_wdat_last     : out std_logic;
      l_linestatus_o_cmd_valid         : in  std_logic;
      l_linestatus_o_cmd_ready         : out std_logic;
      l_linestatus_o_cmd_firstIdx      : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_linestatus_o_cmd_lastIdx       : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_linestatus_o_cmd_ctrl          : in  std_logic_vector(L_LINESTATUS_O_BUS_ADDR_WIDTH*2-1 downto 0);
      l_linestatus_o_cmd_tag           : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_linestatus_o_unl_valid         : out std_logic;
      l_linestatus_o_unl_ready         : in  std_logic;
      l_linestatus_o_unl_tag           : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_sum_qty_valid                  : in  std_logic;
      l_sum_qty_ready                  : out std_logic;
      l_sum_qty_dvalid                 : in  std_logic;
      l_sum_qty_last                   : in  std_logic;
      l_sum_qty                        : in  std_logic_vector(63 downto 0);
      l_sum_qty_bus_wreq_valid         : out std_logic;
      l_sum_qty_bus_wreq_ready         : in  std_logic;
      l_sum_qty_bus_wreq_addr          : out std_logic_vector(L_SUM_QTY_BUS_ADDR_WIDTH-1 downto 0);
      l_sum_qty_bus_wreq_len           : out std_logic_vector(L_SUM_QTY_BUS_LEN_WIDTH-1 downto 0);
      l_sum_qty_bus_wdat_valid         : out std_logic;
      l_sum_qty_bus_wdat_ready         : in  std_logic;
      l_sum_qty_bus_wdat_data          : out std_logic_vector(L_SUM_QTY_BUS_DATA_WIDTH-1 downto 0);
      l_sum_qty_bus_wdat_strobe        : out std_logic_vector(L_SUM_QTY_BUS_DATA_WIDTH/8-1 downto 0);
      l_sum_qty_bus_wdat_last          : out std_logic;
      l_sum_qty_cmd_valid              : in  std_logic;
      l_sum_qty_cmd_ready              : out std_logic;
      l_sum_qty_cmd_firstIdx           : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_sum_qty_cmd_lastIdx            : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_sum_qty_cmd_ctrl               : in  std_logic_vector(L_SUM_QTY_BUS_ADDR_WIDTH-1 downto 0);
      l_sum_qty_cmd_tag                : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_sum_qty_unl_valid              : out std_logic;
      l_sum_qty_unl_ready              : in  std_logic;
      l_sum_qty_unl_tag                : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_sum_base_price_valid           : in  std_logic;
      l_sum_base_price_ready           : out std_logic;
      l_sum_base_price_dvalid          : in  std_logic;
      l_sum_base_price_last            : in  std_logic;
      l_sum_base_price                 : in  std_logic_vector(63 downto 0);
      l_sum_base_price_bus_wreq_valid  : out std_logic;
      l_sum_base_price_bus_wreq_ready  : in  std_logic;
      l_sum_base_price_bus_wreq_addr   : out std_logic_vector(L_SUM_BASE_PRICE_BUS_ADDR_WIDTH-1 downto 0);
      l_sum_base_price_bus_wreq_len    : out std_logic_vector(L_SUM_BASE_PRICE_BUS_LEN_WIDTH-1 downto 0);
      l_sum_base_price_bus_wdat_valid  : out std_logic;
      l_sum_base_price_bus_wdat_ready  : in  std_logic;
      l_sum_base_price_bus_wdat_data   : out std_logic_vector(L_SUM_BASE_PRICE_BUS_DATA_WIDTH-1 downto 0);
      l_sum_base_price_bus_wdat_strobe : out std_logic_vector(L_SUM_BASE_PRICE_BUS_DATA_WIDTH/8-1 downto 0);
      l_sum_base_price_bus_wdat_last   : out std_logic;
      l_sum_base_price_cmd_valid       : in  std_logic;
      l_sum_base_price_cmd_ready       : out std_logic;
      l_sum_base_price_cmd_firstIdx    : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_sum_base_price_cmd_lastIdx     : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_sum_base_price_cmd_ctrl        : in  std_logic_vector(L_SUM_BASE_PRICE_BUS_ADDR_WIDTH-1 downto 0);
      l_sum_base_price_cmd_tag         : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_sum_base_price_unl_valid       : out std_logic;
      l_sum_base_price_unl_ready       : in  std_logic;
      l_sum_base_price_unl_tag         : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_sum_disc_price_valid           : in  std_logic;
      l_sum_disc_price_ready           : out std_logic;
      l_sum_disc_price_dvalid          : in  std_logic;
      l_sum_disc_price_last            : in  std_logic;
      l_sum_disc_price                 : in  std_logic_vector(63 downto 0);
      l_sum_disc_price_bus_wreq_valid  : out std_logic;
      l_sum_disc_price_bus_wreq_ready  : in  std_logic;
      l_sum_disc_price_bus_wreq_addr   : out std_logic_vector(L_SUM_DISC_PRICE_BUS_ADDR_WIDTH-1 downto 0);
      l_sum_disc_price_bus_wreq_len    : out std_logic_vector(L_SUM_DISC_PRICE_BUS_LEN_WIDTH-1 downto 0);
      l_sum_disc_price_bus_wdat_valid  : out std_logic;
      l_sum_disc_price_bus_wdat_ready  : in  std_logic;
      l_sum_disc_price_bus_wdat_data   : out std_logic_vector(L_SUM_DISC_PRICE_BUS_DATA_WIDTH-1 downto 0);
      l_sum_disc_price_bus_wdat_strobe : out std_logic_vector(L_SUM_DISC_PRICE_BUS_DATA_WIDTH/8-1 downto 0);
      l_sum_disc_price_bus_wdat_last   : out std_logic;
      l_sum_disc_price_cmd_valid       : in  std_logic;
      l_sum_disc_price_cmd_ready       : out std_logic;
      l_sum_disc_price_cmd_firstIdx    : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_sum_disc_price_cmd_lastIdx     : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_sum_disc_price_cmd_ctrl        : in  std_logic_vector(L_SUM_DISC_PRICE_BUS_ADDR_WIDTH-1 downto 0);
      l_sum_disc_price_cmd_tag         : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_sum_disc_price_unl_valid       : out std_logic;
      l_sum_disc_price_unl_ready       : in  std_logic;
      l_sum_disc_price_unl_tag         : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_sum_charge_valid               : in  std_logic;
      l_sum_charge_ready               : out std_logic;
      l_sum_charge_dvalid              : in  std_logic;
      l_sum_charge_last                : in  std_logic;
      l_sum_charge                     : in  std_logic_vector(63 downto 0);
      l_sum_charge_bus_wreq_valid      : out std_logic;
      l_sum_charge_bus_wreq_ready      : in  std_logic;
      l_sum_charge_bus_wreq_addr       : out std_logic_vector(L_SUM_CHARGE_BUS_ADDR_WIDTH-1 downto 0);
      l_sum_charge_bus_wreq_len        : out std_logic_vector(L_SUM_CHARGE_BUS_LEN_WIDTH-1 downto 0);
      l_sum_charge_bus_wdat_valid      : out std_logic;
      l_sum_charge_bus_wdat_ready      : in  std_logic;
      l_sum_charge_bus_wdat_data       : out std_logic_vector(L_SUM_CHARGE_BUS_DATA_WIDTH-1 downto 0);
      l_sum_charge_bus_wdat_strobe     : out std_logic_vector(L_SUM_CHARGE_BUS_DATA_WIDTH/8-1 downto 0);
      l_sum_charge_bus_wdat_last       : out std_logic;
      l_sum_charge_cmd_valid           : in  std_logic;
      l_sum_charge_cmd_ready           : out std_logic;
      l_sum_charge_cmd_firstIdx        : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_sum_charge_cmd_lastIdx         : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_sum_charge_cmd_ctrl            : in  std_logic_vector(L_SUM_CHARGE_BUS_ADDR_WIDTH-1 downto 0);
      l_sum_charge_cmd_tag             : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_sum_charge_unl_valid           : out std_logic;
      l_sum_charge_unl_ready           : in  std_logic;
      l_sum_charge_unl_tag             : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_avg_qty_valid                  : in  std_logic;
      l_avg_qty_ready                  : out std_logic;
      l_avg_qty_dvalid                 : in  std_logic;
      l_avg_qty_last                   : in  std_logic;
      l_avg_qty                        : in  std_logic_vector(63 downto 0);
      l_avg_qty_bus_wreq_valid         : out std_logic;
      l_avg_qty_bus_wreq_ready         : in  std_logic;
      l_avg_qty_bus_wreq_addr          : out std_logic_vector(L_AVG_QTY_BUS_ADDR_WIDTH-1 downto 0);
      l_avg_qty_bus_wreq_len           : out std_logic_vector(L_AVG_QTY_BUS_LEN_WIDTH-1 downto 0);
      l_avg_qty_bus_wdat_valid         : out std_logic;
      l_avg_qty_bus_wdat_ready         : in  std_logic;
      l_avg_qty_bus_wdat_data          : out std_logic_vector(L_AVG_QTY_BUS_DATA_WIDTH-1 downto 0);
      l_avg_qty_bus_wdat_strobe        : out std_logic_vector(L_AVG_QTY_BUS_DATA_WIDTH/8-1 downto 0);
      l_avg_qty_bus_wdat_last          : out std_logic;
      l_avg_qty_cmd_valid              : in  std_logic;
      l_avg_qty_cmd_ready              : out std_logic;
      l_avg_qty_cmd_firstIdx           : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_avg_qty_cmd_lastIdx            : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_avg_qty_cmd_ctrl               : in  std_logic_vector(L_AVG_QTY_BUS_ADDR_WIDTH-1 downto 0);
      l_avg_qty_cmd_tag                : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_avg_qty_unl_valid              : out std_logic;
      l_avg_qty_unl_ready              : in  std_logic;
      l_avg_qty_unl_tag                : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_avg_price_valid                : in  std_logic;
      l_avg_price_ready                : out std_logic;
      l_avg_price_dvalid               : in  std_logic;
      l_avg_price_last                 : in  std_logic;
      l_avg_price                      : in  std_logic_vector(63 downto 0);
      l_avg_price_bus_wreq_valid       : out std_logic;
      l_avg_price_bus_wreq_ready       : in  std_logic;
      l_avg_price_bus_wreq_addr        : out std_logic_vector(L_AVG_PRICE_BUS_ADDR_WIDTH-1 downto 0);
      l_avg_price_bus_wreq_len         : out std_logic_vector(L_AVG_PRICE_BUS_LEN_WIDTH-1 downto 0);
      l_avg_price_bus_wdat_valid       : out std_logic;
      l_avg_price_bus_wdat_ready       : in  std_logic;
      l_avg_price_bus_wdat_data        : out std_logic_vector(L_AVG_PRICE_BUS_DATA_WIDTH-1 downto 0);
      l_avg_price_bus_wdat_strobe      : out std_logic_vector(L_AVG_PRICE_BUS_DATA_WIDTH/8-1 downto 0);
      l_avg_price_bus_wdat_last        : out std_logic;
      l_avg_price_cmd_valid            : in  std_logic;
      l_avg_price_cmd_ready            : out std_logic;
      l_avg_price_cmd_firstIdx         : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_avg_price_cmd_lastIdx          : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_avg_price_cmd_ctrl             : in  std_logic_vector(L_AVG_PRICE_BUS_ADDR_WIDTH-1 downto 0);
      l_avg_price_cmd_tag              : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_avg_price_unl_valid            : out std_logic;
      l_avg_price_unl_ready            : in  std_logic;
      l_avg_price_unl_tag              : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_avg_disc_valid                 : in  std_logic;
      l_avg_disc_ready                 : out std_logic;
      l_avg_disc_dvalid                : in  std_logic;
      l_avg_disc_last                  : in  std_logic;
      l_avg_disc                       : in  std_logic_vector(63 downto 0);
      l_avg_disc_bus_wreq_valid        : out std_logic;
      l_avg_disc_bus_wreq_ready        : in  std_logic;
      l_avg_disc_bus_wreq_addr         : out std_logic_vector(L_AVG_DISC_BUS_ADDR_WIDTH-1 downto 0);
      l_avg_disc_bus_wreq_len          : out std_logic_vector(L_AVG_DISC_BUS_LEN_WIDTH-1 downto 0);
      l_avg_disc_bus_wdat_valid        : out std_logic;
      l_avg_disc_bus_wdat_ready        : in  std_logic;
      l_avg_disc_bus_wdat_data         : out std_logic_vector(L_AVG_DISC_BUS_DATA_WIDTH-1 downto 0);
      l_avg_disc_bus_wdat_strobe       : out std_logic_vector(L_AVG_DISC_BUS_DATA_WIDTH/8-1 downto 0);
      l_avg_disc_bus_wdat_last         : out std_logic;
      l_avg_disc_cmd_valid             : in  std_logic;
      l_avg_disc_cmd_ready             : out std_logic;
      l_avg_disc_cmd_firstIdx          : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_avg_disc_cmd_lastIdx           : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_avg_disc_cmd_ctrl              : in  std_logic_vector(L_AVG_DISC_BUS_ADDR_WIDTH-1 downto 0);
      l_avg_disc_cmd_tag               : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_avg_disc_unl_valid             : out std_logic;
      l_avg_disc_unl_ready             : in  std_logic;
      l_avg_disc_unl_tag               : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_count_order_valid              : in  std_logic;
      l_count_order_ready              : out std_logic;
      l_count_order_dvalid             : in  std_logic;
      l_count_order_last               : in  std_logic;
      l_count_order                    : in  std_logic_vector(63 downto 0);
      l_count_order_bus_wreq_valid     : out std_logic;
      l_count_order_bus_wreq_ready     : in  std_logic;
      l_count_order_bus_wreq_addr      : out std_logic_vector(L_COUNT_ORDER_BUS_ADDR_WIDTH-1 downto 0);
      l_count_order_bus_wreq_len       : out std_logic_vector(L_COUNT_ORDER_BUS_LEN_WIDTH-1 downto 0);
      l_count_order_bus_wdat_valid     : out std_logic;
      l_count_order_bus_wdat_ready     : in  std_logic;
      l_count_order_bus_wdat_data      : out std_logic_vector(L_COUNT_ORDER_BUS_DATA_WIDTH-1 downto 0);
      l_count_order_bus_wdat_strobe    : out std_logic_vector(L_COUNT_ORDER_BUS_DATA_WIDTH/8-1 downto 0);
      l_count_order_bus_wdat_last      : out std_logic;
      l_count_order_cmd_valid          : in  std_logic;
      l_count_order_cmd_ready          : out std_logic;
      l_count_order_cmd_firstIdx       : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_count_order_cmd_lastIdx        : in  std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_count_order_cmd_ctrl           : in  std_logic_vector(L_COUNT_ORDER_BUS_ADDR_WIDTH-1 downto 0);
      l_count_order_cmd_tag            : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_count_order_unl_valid          : out std_logic;
      l_count_order_unl_ready          : in  std_logic;
      l_count_order_unl_tag            : out std_logic_vector(TAG_WIDTH-1 downto 0)
    );
  end component;

  signal PriceSummaryWriter_Nucleus_inst_mmio_awvalid                  : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_mmio_awready                  : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_mmio_awaddr                   : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_mmio_wvalid                   : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_mmio_wready                   : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_mmio_wdata                    : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_mmio_wstrb                    : std_logic_vector(3 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_mmio_bvalid                   : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_mmio_bready                   : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_mmio_bresp                    : std_logic_vector(1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_mmio_arvalid                  : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_mmio_arready                  : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_mmio_araddr                   : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_mmio_rvalid                   : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_mmio_rready                   : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_mmio_rdata                    : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_mmio_rresp                    : std_logic_vector(1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_valid          : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_ready          : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_dvalid         : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_last           : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_length         : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_count          : std_logic_vector(0 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_valid    : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_ready    : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_dvalid   : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_last     : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars          : std_logic_vector(7 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_count    : std_logic_vector(0 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_valid          : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_ready          : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_dvalid         : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_last           : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_length         : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_count          : std_logic_vector(0 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_valid    : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_ready    : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_dvalid   : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_last     : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars          : std_logic_vector(7 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_count    : std_logic_vector(0 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_sum_qty_valid               : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_qty_ready               : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_qty_dvalid              : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_qty_last                : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_qty                     : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_sum_base_price_valid        : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_base_price_ready        : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_base_price_dvalid       : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_base_price_last         : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_base_price              : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_valid        : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_ready        : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_dvalid       : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_last         : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_disc_price              : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_sum_charge_valid            : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_charge_ready            : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_charge_dvalid           : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_charge_last             : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_charge                  : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_avg_qty_valid               : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_qty_ready               : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_qty_dvalid              : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_qty_last                : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_qty                     : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_avg_price_valid             : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_price_ready             : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_price_dvalid            : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_price_last              : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_price                   : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_avg_disc_valid              : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_disc_ready              : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_disc_dvalid             : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_disc_last               : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_disc                    : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_count_order_valid           : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_count_order_ready           : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_count_order_dvalid          : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_count_order_last            : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_count_order                 : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_unl_valid      : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_unl_ready      : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_unl_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_unl_valid      : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_unl_ready      : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_unl_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_sum_qty_unl_valid           : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_qty_unl_ready           : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_qty_unl_tag             : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_sum_base_price_unl_valid    : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_base_price_unl_ready    : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_base_price_unl_tag      : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_unl_valid    : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_unl_ready    : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_unl_tag      : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_sum_charge_unl_valid        : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_charge_unl_ready        : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_charge_unl_tag          : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_avg_qty_unl_valid           : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_qty_unl_ready           : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_qty_unl_tag             : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_avg_price_unl_valid         : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_price_unl_ready         : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_price_unl_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_avg_disc_unl_valid          : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_disc_unl_ready          : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_disc_unl_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_count_order_unl_valid       : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_count_order_unl_ready       : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_count_order_unl_tag         : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_valid      : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_ready      : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_firstIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_lastIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_ctrl       : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_valid      : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_ready      : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_firstIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_lastIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_ctrl       : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_tag        : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_valid           : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_ready           : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_firstIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_lastIdx         : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_ctrl            : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_tag             : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_valid    : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_ready    : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_firstIdx : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_lastIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_ctrl     : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_tag      : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_valid    : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_ready    : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_firstIdx : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_lastIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_ctrl     : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_tag      : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_valid        : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_ready        : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_firstIdx     : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_lastIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_ctrl         : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_tag          : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_valid           : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_ready           : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_firstIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_lastIdx         : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_ctrl            : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_tag             : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_valid         : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_ready         : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_ctrl          : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_valid          : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_ready          : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_ctrl           : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_valid       : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_ready       : std_logic;
  signal PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_firstIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_lastIdx     : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_ctrl        : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_tag         : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_l_inst_l_returnflag_o_valid                : std_logic;
  signal PriceSummaryWriter_l_inst_l_returnflag_o_ready                : std_logic;
  signal PriceSummaryWriter_l_inst_l_returnflag_o_dvalid               : std_logic;
  signal PriceSummaryWriter_l_inst_l_returnflag_o_last                 : std_logic;
  signal PriceSummaryWriter_l_inst_l_returnflag_o_length               : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_l_inst_l_returnflag_o_count                : std_logic_vector(0 downto 0);
  signal PriceSummaryWriter_l_inst_l_returnflag_o_chars_valid          : std_logic;
  signal PriceSummaryWriter_l_inst_l_returnflag_o_chars_ready          : std_logic;
  signal PriceSummaryWriter_l_inst_l_returnflag_o_chars_dvalid         : std_logic;
  signal PriceSummaryWriter_l_inst_l_returnflag_o_chars_last           : std_logic;
  signal PriceSummaryWriter_l_inst_l_returnflag_o_chars                : std_logic_vector(7 downto 0);
  signal PriceSummaryWriter_l_inst_l_returnflag_o_chars_count          : std_logic_vector(0 downto 0);

  signal PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_valid       : std_logic;
  signal PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_ready       : std_logic;
  signal PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_addr        : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_len         : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_valid       : std_logic;
  signal PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_ready       : std_logic;
  signal PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_data        : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_strobe      : std_logic_vector(BUS_DATA_WIDTH/8-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_last        : std_logic;

  signal PriceSummaryWriter_l_inst_l_returnflag_o_cmd_valid            : std_logic;
  signal PriceSummaryWriter_l_inst_l_returnflag_o_cmd_ready            : std_logic;
  signal PriceSummaryWriter_l_inst_l_returnflag_o_cmd_firstIdx         : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_returnflag_o_cmd_lastIdx          : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_returnflag_o_cmd_ctrl             : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_returnflag_o_cmd_tag              : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_l_inst_l_returnflag_o_unl_valid            : std_logic;
  signal PriceSummaryWriter_l_inst_l_returnflag_o_unl_ready            : std_logic;
  signal PriceSummaryWriter_l_inst_l_returnflag_o_unl_tag              : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_l_inst_l_linestatus_o_valid                : std_logic;
  signal PriceSummaryWriter_l_inst_l_linestatus_o_ready                : std_logic;
  signal PriceSummaryWriter_l_inst_l_linestatus_o_dvalid               : std_logic;
  signal PriceSummaryWriter_l_inst_l_linestatus_o_last                 : std_logic;
  signal PriceSummaryWriter_l_inst_l_linestatus_o_length               : std_logic_vector(31 downto 0);
  signal PriceSummaryWriter_l_inst_l_linestatus_o_count                : std_logic_vector(0 downto 0);
  signal PriceSummaryWriter_l_inst_l_linestatus_o_chars_valid          : std_logic;
  signal PriceSummaryWriter_l_inst_l_linestatus_o_chars_ready          : std_logic;
  signal PriceSummaryWriter_l_inst_l_linestatus_o_chars_dvalid         : std_logic;
  signal PriceSummaryWriter_l_inst_l_linestatus_o_chars_last           : std_logic;
  signal PriceSummaryWriter_l_inst_l_linestatus_o_chars                : std_logic_vector(7 downto 0);
  signal PriceSummaryWriter_l_inst_l_linestatus_o_chars_count          : std_logic_vector(0 downto 0);

  signal PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_valid       : std_logic;
  signal PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_ready       : std_logic;
  signal PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_addr        : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_len         : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_valid       : std_logic;
  signal PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_ready       : std_logic;
  signal PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_data        : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_strobe      : std_logic_vector(BUS_DATA_WIDTH/8-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_last        : std_logic;

  signal PriceSummaryWriter_l_inst_l_linestatus_o_cmd_valid            : std_logic;
  signal PriceSummaryWriter_l_inst_l_linestatus_o_cmd_ready            : std_logic;
  signal PriceSummaryWriter_l_inst_l_linestatus_o_cmd_firstIdx         : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_linestatus_o_cmd_lastIdx          : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_linestatus_o_cmd_ctrl             : std_logic_vector(BUS_ADDR_WIDTH*2-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_linestatus_o_cmd_tag              : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_l_inst_l_linestatus_o_unl_valid            : std_logic;
  signal PriceSummaryWriter_l_inst_l_linestatus_o_unl_ready            : std_logic;
  signal PriceSummaryWriter_l_inst_l_linestatus_o_unl_tag              : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_l_inst_l_sum_qty_valid                     : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_qty_ready                     : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_qty_dvalid                    : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_qty_last                      : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_qty                           : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_valid            : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_ready            : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_addr             : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_len              : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_valid            : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_ready            : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_data             : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_strobe           : std_logic_vector(BUS_DATA_WIDTH/8-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_last             : std_logic;

  signal PriceSummaryWriter_l_inst_l_sum_qty_cmd_valid                 : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_qty_cmd_ready                 : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_qty_cmd_firstIdx              : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_qty_cmd_lastIdx               : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_qty_cmd_ctrl                  : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_qty_cmd_tag                   : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_l_inst_l_sum_qty_unl_valid                 : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_qty_unl_ready                 : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_qty_unl_tag                   : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_l_inst_l_sum_base_price_valid              : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_base_price_ready              : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_base_price_dvalid             : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_base_price_last               : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_base_price                    : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_valid     : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_ready     : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_addr      : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_len       : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_valid     : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_ready     : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_data      : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_strobe    : std_logic_vector(BUS_DATA_WIDTH/8-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_last      : std_logic;

  signal PriceSummaryWriter_l_inst_l_sum_base_price_cmd_valid          : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_base_price_cmd_ready          : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_base_price_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_base_price_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_base_price_cmd_ctrl           : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_base_price_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_l_inst_l_sum_base_price_unl_valid          : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_base_price_unl_ready          : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_base_price_unl_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_l_inst_l_sum_disc_price_valid              : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_ready              : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_dvalid             : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_last               : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_disc_price                    : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_valid     : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_ready     : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_addr      : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_len       : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_valid     : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_ready     : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_data      : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_strobe    : std_logic_vector(BUS_DATA_WIDTH/8-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_last      : std_logic;

  signal PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_valid          : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_ready          : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_ctrl           : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_l_inst_l_sum_disc_price_unl_valid          : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_unl_ready          : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_disc_price_unl_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_l_inst_l_sum_charge_valid                  : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_charge_ready                  : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_charge_dvalid                 : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_charge_last                   : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_charge                        : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_valid         : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_ready         : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_addr          : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_len           : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_valid         : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_ready         : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_data          : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_strobe        : std_logic_vector(BUS_DATA_WIDTH/8-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_last          : std_logic;

  signal PriceSummaryWriter_l_inst_l_sum_charge_cmd_valid              : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_charge_cmd_ready              : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_charge_cmd_firstIdx           : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_charge_cmd_lastIdx            : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_charge_cmd_ctrl               : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_sum_charge_cmd_tag                : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_l_inst_l_sum_charge_unl_valid              : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_charge_unl_ready              : std_logic;
  signal PriceSummaryWriter_l_inst_l_sum_charge_unl_tag                : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_l_inst_l_avg_qty_valid                     : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_qty_ready                     : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_qty_dvalid                    : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_qty_last                      : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_qty                           : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_valid            : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_ready            : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_addr             : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_len              : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_valid            : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_ready            : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_data             : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_strobe           : std_logic_vector(BUS_DATA_WIDTH/8-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_last             : std_logic;

  signal PriceSummaryWriter_l_inst_l_avg_qty_cmd_valid                 : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_qty_cmd_ready                 : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_qty_cmd_firstIdx              : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_qty_cmd_lastIdx               : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_qty_cmd_ctrl                  : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_qty_cmd_tag                   : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_l_inst_l_avg_qty_unl_valid                 : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_qty_unl_ready                 : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_qty_unl_tag                   : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_l_inst_l_avg_price_valid                   : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_price_ready                   : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_price_dvalid                  : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_price_last                    : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_price                         : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_valid          : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_ready          : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_addr           : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_len            : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_valid          : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_ready          : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_data           : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_strobe         : std_logic_vector(BUS_DATA_WIDTH/8-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_last           : std_logic;

  signal PriceSummaryWriter_l_inst_l_avg_price_cmd_valid               : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_price_cmd_ready               : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_price_cmd_firstIdx            : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_price_cmd_lastIdx             : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_price_cmd_ctrl                : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_price_cmd_tag                 : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_l_inst_l_avg_price_unl_valid               : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_price_unl_ready               : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_price_unl_tag                 : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_l_inst_l_avg_disc_valid                    : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_disc_ready                    : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_disc_dvalid                   : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_disc_last                     : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_disc                          : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_valid           : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_ready           : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_addr            : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_len             : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_valid           : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_ready           : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_data            : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_strobe          : std_logic_vector(BUS_DATA_WIDTH/8-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_last            : std_logic;

  signal PriceSummaryWriter_l_inst_l_avg_disc_cmd_valid                : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_disc_cmd_ready                : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_disc_cmd_firstIdx             : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_disc_cmd_lastIdx              : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_disc_cmd_ctrl                 : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_avg_disc_cmd_tag                  : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_l_inst_l_avg_disc_unl_valid                : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_disc_unl_ready                : std_logic;
  signal PriceSummaryWriter_l_inst_l_avg_disc_unl_tag                  : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_l_inst_l_count_order_valid                 : std_logic;
  signal PriceSummaryWriter_l_inst_l_count_order_ready                 : std_logic;
  signal PriceSummaryWriter_l_inst_l_count_order_dvalid                : std_logic;
  signal PriceSummaryWriter_l_inst_l_count_order_last                  : std_logic;
  signal PriceSummaryWriter_l_inst_l_count_order                       : std_logic_vector(63 downto 0);

  signal PriceSummaryWriter_l_inst_l_count_order_bus_wreq_valid        : std_logic;
  signal PriceSummaryWriter_l_inst_l_count_order_bus_wreq_ready        : std_logic;
  signal PriceSummaryWriter_l_inst_l_count_order_bus_wreq_addr         : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_count_order_bus_wreq_len          : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_count_order_bus_wdat_valid        : std_logic;
  signal PriceSummaryWriter_l_inst_l_count_order_bus_wdat_ready        : std_logic;
  signal PriceSummaryWriter_l_inst_l_count_order_bus_wdat_data         : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_count_order_bus_wdat_strobe       : std_logic_vector(BUS_DATA_WIDTH/8-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_count_order_bus_wdat_last         : std_logic;

  signal PriceSummaryWriter_l_inst_l_count_order_cmd_valid             : std_logic;
  signal PriceSummaryWriter_l_inst_l_count_order_cmd_ready             : std_logic;
  signal PriceSummaryWriter_l_inst_l_count_order_cmd_firstIdx          : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_count_order_cmd_lastIdx           : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_count_order_cmd_ctrl              : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal PriceSummaryWriter_l_inst_l_count_order_cmd_tag               : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal PriceSummaryWriter_l_inst_l_count_order_unl_valid             : std_logic;
  signal PriceSummaryWriter_l_inst_l_count_order_unl_ready             : std_logic;
  signal PriceSummaryWriter_l_inst_l_count_order_unl_tag               : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal WRAW64DW512LW8BS1BM16_inst_mst_wreq_valid                     : std_logic;
  signal WRAW64DW512LW8BS1BM16_inst_mst_wreq_ready                     : std_logic;
  signal WRAW64DW512LW8BS1BM16_inst_mst_wreq_addr                      : std_logic_vector(BUS_ADDR_WIDTH-1 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_mst_wreq_len                       : std_logic_vector(BUS_LEN_WIDTH-1 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_mst_wdat_valid                     : std_logic;
  signal WRAW64DW512LW8BS1BM16_inst_mst_wdat_ready                     : std_logic;
  signal WRAW64DW512LW8BS1BM16_inst_mst_wdat_data                      : std_logic_vector(BUS_DATA_WIDTH-1 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_mst_wdat_strobe                    : std_logic_vector(BUS_DATA_WIDTH/8-1 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_mst_wdat_last                      : std_logic;

  signal WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid  : std_logic_vector(9 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready  : std_logic_vector(9 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr   : std_logic_vector(10*BUS_ADDR_WIDTH-1 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len    : std_logic_vector(10*BUS_LEN_WIDTH-1 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid  : std_logic_vector(9 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready  : std_logic_vector(9 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data   : std_logic_vector(10*BUS_DATA_WIDTH-1 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe : std_logic_vector(10*BUS_DATA_WIDTH/8-1 downto 0);
  signal WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last   : std_logic_vector(9 downto 0);

begin
  PriceSummaryWriter_Nucleus_inst : PriceSummaryWriter_Nucleus
    generic map (
      INDEX_WIDTH                     => INDEX_WIDTH,
      TAG_WIDTH                       => TAG_WIDTH,
      L_RETURNFLAG_O_BUS_ADDR_WIDTH   => BUS_ADDR_WIDTH,
      L_LINESTATUS_O_BUS_ADDR_WIDTH   => BUS_ADDR_WIDTH,
      L_SUM_QTY_BUS_ADDR_WIDTH        => BUS_ADDR_WIDTH,
      L_SUM_BASE_PRICE_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
      L_SUM_DISC_PRICE_BUS_ADDR_WIDTH => BUS_ADDR_WIDTH,
      L_SUM_CHARGE_BUS_ADDR_WIDTH     => BUS_ADDR_WIDTH,
      L_AVG_QTY_BUS_ADDR_WIDTH        => BUS_ADDR_WIDTH,
      L_AVG_PRICE_BUS_ADDR_WIDTH      => BUS_ADDR_WIDTH,
      L_AVG_DISC_BUS_ADDR_WIDTH       => BUS_ADDR_WIDTH,
      L_COUNT_ORDER_BUS_ADDR_WIDTH    => BUS_ADDR_WIDTH
    )
    port map (
      kcd_clk                       => kcd_clk,
      kcd_reset                     => kcd_reset,
      mmio_awvalid                  => PriceSummaryWriter_Nucleus_inst_mmio_awvalid,
      mmio_awready                  => PriceSummaryWriter_Nucleus_inst_mmio_awready,
      mmio_awaddr                   => PriceSummaryWriter_Nucleus_inst_mmio_awaddr,
      mmio_wvalid                   => PriceSummaryWriter_Nucleus_inst_mmio_wvalid,
      mmio_wready                   => PriceSummaryWriter_Nucleus_inst_mmio_wready,
      mmio_wdata                    => PriceSummaryWriter_Nucleus_inst_mmio_wdata,
      mmio_wstrb                    => PriceSummaryWriter_Nucleus_inst_mmio_wstrb,
      mmio_bvalid                   => PriceSummaryWriter_Nucleus_inst_mmio_bvalid,
      mmio_bready                   => PriceSummaryWriter_Nucleus_inst_mmio_bready,
      mmio_bresp                    => PriceSummaryWriter_Nucleus_inst_mmio_bresp,
      mmio_arvalid                  => PriceSummaryWriter_Nucleus_inst_mmio_arvalid,
      mmio_arready                  => PriceSummaryWriter_Nucleus_inst_mmio_arready,
      mmio_araddr                   => PriceSummaryWriter_Nucleus_inst_mmio_araddr,
      mmio_rvalid                   => PriceSummaryWriter_Nucleus_inst_mmio_rvalid,
      mmio_rready                   => PriceSummaryWriter_Nucleus_inst_mmio_rready,
      mmio_rdata                    => PriceSummaryWriter_Nucleus_inst_mmio_rdata,
      mmio_rresp                    => PriceSummaryWriter_Nucleus_inst_mmio_rresp,
      l_returnflag_o_valid          => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_valid,
      l_returnflag_o_ready          => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_ready,
      l_returnflag_o_dvalid         => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_dvalid,
      l_returnflag_o_last           => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_last,
      l_returnflag_o_length         => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_length,
      l_returnflag_o_count          => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_count,
      l_returnflag_o_chars_valid    => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_valid,
      l_returnflag_o_chars_ready    => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_ready,
      l_returnflag_o_chars_dvalid   => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_dvalid,
      l_returnflag_o_chars_last     => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_last,
      l_returnflag_o_chars          => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars,
      l_returnflag_o_chars_count    => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_count,
      l_linestatus_o_valid          => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_valid,
      l_linestatus_o_ready          => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_ready,
      l_linestatus_o_dvalid         => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_dvalid,
      l_linestatus_o_last           => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_last,
      l_linestatus_o_length         => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_length,
      l_linestatus_o_count          => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_count,
      l_linestatus_o_chars_valid    => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_valid,
      l_linestatus_o_chars_ready    => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_ready,
      l_linestatus_o_chars_dvalid   => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_dvalid,
      l_linestatus_o_chars_last     => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_last,
      l_linestatus_o_chars          => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars,
      l_linestatus_o_chars_count    => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_count,
      l_sum_qty_valid               => PriceSummaryWriter_Nucleus_inst_l_sum_qty_valid,
      l_sum_qty_ready               => PriceSummaryWriter_Nucleus_inst_l_sum_qty_ready,
      l_sum_qty_dvalid              => PriceSummaryWriter_Nucleus_inst_l_sum_qty_dvalid,
      l_sum_qty_last                => PriceSummaryWriter_Nucleus_inst_l_sum_qty_last,
      l_sum_qty                     => PriceSummaryWriter_Nucleus_inst_l_sum_qty,
      l_sum_base_price_valid        => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_valid,
      l_sum_base_price_ready        => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_ready,
      l_sum_base_price_dvalid       => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_dvalid,
      l_sum_base_price_last         => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_last,
      l_sum_base_price              => PriceSummaryWriter_Nucleus_inst_l_sum_base_price,
      l_sum_disc_price_valid        => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_valid,
      l_sum_disc_price_ready        => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_ready,
      l_sum_disc_price_dvalid       => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_dvalid,
      l_sum_disc_price_last         => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_last,
      l_sum_disc_price              => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price,
      l_sum_charge_valid            => PriceSummaryWriter_Nucleus_inst_l_sum_charge_valid,
      l_sum_charge_ready            => PriceSummaryWriter_Nucleus_inst_l_sum_charge_ready,
      l_sum_charge_dvalid           => PriceSummaryWriter_Nucleus_inst_l_sum_charge_dvalid,
      l_sum_charge_last             => PriceSummaryWriter_Nucleus_inst_l_sum_charge_last,
      l_sum_charge                  => PriceSummaryWriter_Nucleus_inst_l_sum_charge,
      l_avg_qty_valid               => PriceSummaryWriter_Nucleus_inst_l_avg_qty_valid,
      l_avg_qty_ready               => PriceSummaryWriter_Nucleus_inst_l_avg_qty_ready,
      l_avg_qty_dvalid              => PriceSummaryWriter_Nucleus_inst_l_avg_qty_dvalid,
      l_avg_qty_last                => PriceSummaryWriter_Nucleus_inst_l_avg_qty_last,
      l_avg_qty                     => PriceSummaryWriter_Nucleus_inst_l_avg_qty,
      l_avg_price_valid             => PriceSummaryWriter_Nucleus_inst_l_avg_price_valid,
      l_avg_price_ready             => PriceSummaryWriter_Nucleus_inst_l_avg_price_ready,
      l_avg_price_dvalid            => PriceSummaryWriter_Nucleus_inst_l_avg_price_dvalid,
      l_avg_price_last              => PriceSummaryWriter_Nucleus_inst_l_avg_price_last,
      l_avg_price                   => PriceSummaryWriter_Nucleus_inst_l_avg_price,
      l_avg_disc_valid              => PriceSummaryWriter_Nucleus_inst_l_avg_disc_valid,
      l_avg_disc_ready              => PriceSummaryWriter_Nucleus_inst_l_avg_disc_ready,
      l_avg_disc_dvalid             => PriceSummaryWriter_Nucleus_inst_l_avg_disc_dvalid,
      l_avg_disc_last               => PriceSummaryWriter_Nucleus_inst_l_avg_disc_last,
      l_avg_disc                    => PriceSummaryWriter_Nucleus_inst_l_avg_disc,
      l_count_order_valid           => PriceSummaryWriter_Nucleus_inst_l_count_order_valid,
      l_count_order_ready           => PriceSummaryWriter_Nucleus_inst_l_count_order_ready,
      l_count_order_dvalid          => PriceSummaryWriter_Nucleus_inst_l_count_order_dvalid,
      l_count_order_last            => PriceSummaryWriter_Nucleus_inst_l_count_order_last,
      l_count_order                 => PriceSummaryWriter_Nucleus_inst_l_count_order,
      l_returnflag_o_unl_valid      => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_unl_valid,
      l_returnflag_o_unl_ready      => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_unl_ready,
      l_returnflag_o_unl_tag        => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_unl_tag,
      l_linestatus_o_unl_valid      => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_unl_valid,
      l_linestatus_o_unl_ready      => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_unl_ready,
      l_linestatus_o_unl_tag        => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_unl_tag,
      l_sum_qty_unl_valid           => PriceSummaryWriter_Nucleus_inst_l_sum_qty_unl_valid,
      l_sum_qty_unl_ready           => PriceSummaryWriter_Nucleus_inst_l_sum_qty_unl_ready,
      l_sum_qty_unl_tag             => PriceSummaryWriter_Nucleus_inst_l_sum_qty_unl_tag,
      l_sum_base_price_unl_valid    => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_unl_valid,
      l_sum_base_price_unl_ready    => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_unl_ready,
      l_sum_base_price_unl_tag      => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_unl_tag,
      l_sum_disc_price_unl_valid    => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_unl_valid,
      l_sum_disc_price_unl_ready    => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_unl_ready,
      l_sum_disc_price_unl_tag      => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_unl_tag,
      l_sum_charge_unl_valid        => PriceSummaryWriter_Nucleus_inst_l_sum_charge_unl_valid,
      l_sum_charge_unl_ready        => PriceSummaryWriter_Nucleus_inst_l_sum_charge_unl_ready,
      l_sum_charge_unl_tag          => PriceSummaryWriter_Nucleus_inst_l_sum_charge_unl_tag,
      l_avg_qty_unl_valid           => PriceSummaryWriter_Nucleus_inst_l_avg_qty_unl_valid,
      l_avg_qty_unl_ready           => PriceSummaryWriter_Nucleus_inst_l_avg_qty_unl_ready,
      l_avg_qty_unl_tag             => PriceSummaryWriter_Nucleus_inst_l_avg_qty_unl_tag,
      l_avg_price_unl_valid         => PriceSummaryWriter_Nucleus_inst_l_avg_price_unl_valid,
      l_avg_price_unl_ready         => PriceSummaryWriter_Nucleus_inst_l_avg_price_unl_ready,
      l_avg_price_unl_tag           => PriceSummaryWriter_Nucleus_inst_l_avg_price_unl_tag,
      l_avg_disc_unl_valid          => PriceSummaryWriter_Nucleus_inst_l_avg_disc_unl_valid,
      l_avg_disc_unl_ready          => PriceSummaryWriter_Nucleus_inst_l_avg_disc_unl_ready,
      l_avg_disc_unl_tag            => PriceSummaryWriter_Nucleus_inst_l_avg_disc_unl_tag,
      l_count_order_unl_valid       => PriceSummaryWriter_Nucleus_inst_l_count_order_unl_valid,
      l_count_order_unl_ready       => PriceSummaryWriter_Nucleus_inst_l_count_order_unl_ready,
      l_count_order_unl_tag         => PriceSummaryWriter_Nucleus_inst_l_count_order_unl_tag,
      l_returnflag_o_cmd_valid      => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_valid,
      l_returnflag_o_cmd_ready      => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_ready,
      l_returnflag_o_cmd_firstIdx   => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_firstIdx,
      l_returnflag_o_cmd_lastIdx    => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_lastIdx,
      l_returnflag_o_cmd_ctrl       => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_ctrl,
      l_returnflag_o_cmd_tag        => PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_tag,
      l_linestatus_o_cmd_valid      => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_valid,
      l_linestatus_o_cmd_ready      => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_ready,
      l_linestatus_o_cmd_firstIdx   => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_firstIdx,
      l_linestatus_o_cmd_lastIdx    => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_lastIdx,
      l_linestatus_o_cmd_ctrl       => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_ctrl,
      l_linestatus_o_cmd_tag        => PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_tag,
      l_sum_qty_cmd_valid           => PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_valid,
      l_sum_qty_cmd_ready           => PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_ready,
      l_sum_qty_cmd_firstIdx        => PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_firstIdx,
      l_sum_qty_cmd_lastIdx         => PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_lastIdx,
      l_sum_qty_cmd_ctrl            => PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_ctrl,
      l_sum_qty_cmd_tag             => PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_tag,
      l_sum_base_price_cmd_valid    => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_valid,
      l_sum_base_price_cmd_ready    => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_ready,
      l_sum_base_price_cmd_firstIdx => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_firstIdx,
      l_sum_base_price_cmd_lastIdx  => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_lastIdx,
      l_sum_base_price_cmd_ctrl     => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_ctrl,
      l_sum_base_price_cmd_tag      => PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_tag,
      l_sum_disc_price_cmd_valid    => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_valid,
      l_sum_disc_price_cmd_ready    => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_ready,
      l_sum_disc_price_cmd_firstIdx => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_firstIdx,
      l_sum_disc_price_cmd_lastIdx  => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_lastIdx,
      l_sum_disc_price_cmd_ctrl     => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_ctrl,
      l_sum_disc_price_cmd_tag      => PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_tag,
      l_sum_charge_cmd_valid        => PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_valid,
      l_sum_charge_cmd_ready        => PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_ready,
      l_sum_charge_cmd_firstIdx     => PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_firstIdx,
      l_sum_charge_cmd_lastIdx      => PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_lastIdx,
      l_sum_charge_cmd_ctrl         => PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_ctrl,
      l_sum_charge_cmd_tag          => PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_tag,
      l_avg_qty_cmd_valid           => PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_valid,
      l_avg_qty_cmd_ready           => PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_ready,
      l_avg_qty_cmd_firstIdx        => PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_firstIdx,
      l_avg_qty_cmd_lastIdx         => PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_lastIdx,
      l_avg_qty_cmd_ctrl            => PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_ctrl,
      l_avg_qty_cmd_tag             => PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_tag,
      l_avg_price_cmd_valid         => PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_valid,
      l_avg_price_cmd_ready         => PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_ready,
      l_avg_price_cmd_firstIdx      => PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_firstIdx,
      l_avg_price_cmd_lastIdx       => PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_lastIdx,
      l_avg_price_cmd_ctrl          => PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_ctrl,
      l_avg_price_cmd_tag           => PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_tag,
      l_avg_disc_cmd_valid          => PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_valid,
      l_avg_disc_cmd_ready          => PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_ready,
      l_avg_disc_cmd_firstIdx       => PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_firstIdx,
      l_avg_disc_cmd_lastIdx        => PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_lastIdx,
      l_avg_disc_cmd_ctrl           => PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_ctrl,
      l_avg_disc_cmd_tag            => PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_tag,
      l_count_order_cmd_valid       => PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_valid,
      l_count_order_cmd_ready       => PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_ready,
      l_count_order_cmd_firstIdx    => PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_firstIdx,
      l_count_order_cmd_lastIdx     => PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_lastIdx,
      l_count_order_cmd_ctrl        => PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_ctrl,
      l_count_order_cmd_tag         => PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_tag
    );

  PriceSummaryWriter_l_inst : PriceSummaryWriter_l
    generic map (
      INDEX_WIDTH                         => INDEX_WIDTH,
      TAG_WIDTH                           => TAG_WIDTH,
      L_RETURNFLAG_O_BUS_ADDR_WIDTH       => BUS_ADDR_WIDTH,
      L_RETURNFLAG_O_BUS_DATA_WIDTH       => BUS_DATA_WIDTH,
      L_RETURNFLAG_O_BUS_LEN_WIDTH        => BUS_LEN_WIDTH,
      L_RETURNFLAG_O_BUS_BURST_STEP_LEN   => BUS_BURST_STEP_LEN,
      L_RETURNFLAG_O_BUS_BURST_MAX_LEN    => BUS_BURST_MAX_LEN,
      L_LINESTATUS_O_BUS_ADDR_WIDTH       => BUS_ADDR_WIDTH,
      L_LINESTATUS_O_BUS_DATA_WIDTH       => BUS_DATA_WIDTH,
      L_LINESTATUS_O_BUS_LEN_WIDTH        => BUS_LEN_WIDTH,
      L_LINESTATUS_O_BUS_BURST_STEP_LEN   => BUS_BURST_STEP_LEN,
      L_LINESTATUS_O_BUS_BURST_MAX_LEN    => BUS_BURST_MAX_LEN,
      L_SUM_QTY_BUS_ADDR_WIDTH            => BUS_ADDR_WIDTH,
      L_SUM_QTY_BUS_DATA_WIDTH            => BUS_DATA_WIDTH,
      L_SUM_QTY_BUS_LEN_WIDTH             => BUS_LEN_WIDTH,
      L_SUM_QTY_BUS_BURST_STEP_LEN        => BUS_BURST_STEP_LEN,
      L_SUM_QTY_BUS_BURST_MAX_LEN         => BUS_BURST_MAX_LEN,
      L_SUM_BASE_PRICE_BUS_ADDR_WIDTH     => BUS_ADDR_WIDTH,
      L_SUM_BASE_PRICE_BUS_DATA_WIDTH     => BUS_DATA_WIDTH,
      L_SUM_BASE_PRICE_BUS_LEN_WIDTH      => BUS_LEN_WIDTH,
      L_SUM_BASE_PRICE_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
      L_SUM_BASE_PRICE_BUS_BURST_MAX_LEN  => BUS_BURST_MAX_LEN,
      L_SUM_DISC_PRICE_BUS_ADDR_WIDTH     => BUS_ADDR_WIDTH,
      L_SUM_DISC_PRICE_BUS_DATA_WIDTH     => BUS_DATA_WIDTH,
      L_SUM_DISC_PRICE_BUS_LEN_WIDTH      => BUS_LEN_WIDTH,
      L_SUM_DISC_PRICE_BUS_BURST_STEP_LEN => BUS_BURST_STEP_LEN,
      L_SUM_DISC_PRICE_BUS_BURST_MAX_LEN  => BUS_BURST_MAX_LEN,
      L_SUM_CHARGE_BUS_ADDR_WIDTH         => BUS_ADDR_WIDTH,
      L_SUM_CHARGE_BUS_DATA_WIDTH         => BUS_DATA_WIDTH,
      L_SUM_CHARGE_BUS_LEN_WIDTH          => BUS_LEN_WIDTH,
      L_SUM_CHARGE_BUS_BURST_STEP_LEN     => BUS_BURST_STEP_LEN,
      L_SUM_CHARGE_BUS_BURST_MAX_LEN      => BUS_BURST_MAX_LEN,
      L_AVG_QTY_BUS_ADDR_WIDTH            => BUS_ADDR_WIDTH,
      L_AVG_QTY_BUS_DATA_WIDTH            => BUS_DATA_WIDTH,
      L_AVG_QTY_BUS_LEN_WIDTH             => BUS_LEN_WIDTH,
      L_AVG_QTY_BUS_BURST_STEP_LEN        => BUS_BURST_STEP_LEN,
      L_AVG_QTY_BUS_BURST_MAX_LEN         => BUS_BURST_MAX_LEN,
      L_AVG_PRICE_BUS_ADDR_WIDTH          => BUS_ADDR_WIDTH,
      L_AVG_PRICE_BUS_DATA_WIDTH          => BUS_DATA_WIDTH,
      L_AVG_PRICE_BUS_LEN_WIDTH           => BUS_LEN_WIDTH,
      L_AVG_PRICE_BUS_BURST_STEP_LEN      => BUS_BURST_STEP_LEN,
      L_AVG_PRICE_BUS_BURST_MAX_LEN       => BUS_BURST_MAX_LEN,
      L_AVG_DISC_BUS_ADDR_WIDTH           => BUS_ADDR_WIDTH,
      L_AVG_DISC_BUS_DATA_WIDTH           => BUS_DATA_WIDTH,
      L_AVG_DISC_BUS_LEN_WIDTH            => BUS_LEN_WIDTH,
      L_AVG_DISC_BUS_BURST_STEP_LEN       => BUS_BURST_STEP_LEN,
      L_AVG_DISC_BUS_BURST_MAX_LEN        => BUS_BURST_MAX_LEN,
      L_COUNT_ORDER_BUS_ADDR_WIDTH        => BUS_ADDR_WIDTH,
      L_COUNT_ORDER_BUS_DATA_WIDTH        => BUS_DATA_WIDTH,
      L_COUNT_ORDER_BUS_LEN_WIDTH         => BUS_LEN_WIDTH,
      L_COUNT_ORDER_BUS_BURST_STEP_LEN    => BUS_BURST_STEP_LEN,
      L_COUNT_ORDER_BUS_BURST_MAX_LEN     => BUS_BURST_MAX_LEN
    )
    port map (
      bcd_clk                          => bcd_clk,
      bcd_reset                        => bcd_reset,
      kcd_clk                          => kcd_clk,
      kcd_reset                        => kcd_reset,
      l_returnflag_o_valid             => PriceSummaryWriter_l_inst_l_returnflag_o_valid,
      l_returnflag_o_ready             => PriceSummaryWriter_l_inst_l_returnflag_o_ready,
      l_returnflag_o_dvalid            => PriceSummaryWriter_l_inst_l_returnflag_o_dvalid,
      l_returnflag_o_last              => PriceSummaryWriter_l_inst_l_returnflag_o_last,
      l_returnflag_o_length            => PriceSummaryWriter_l_inst_l_returnflag_o_length,
      l_returnflag_o_count             => PriceSummaryWriter_l_inst_l_returnflag_o_count,
      l_returnflag_o_chars_valid       => PriceSummaryWriter_l_inst_l_returnflag_o_chars_valid,
      l_returnflag_o_chars_ready       => PriceSummaryWriter_l_inst_l_returnflag_o_chars_ready,
      l_returnflag_o_chars_dvalid      => PriceSummaryWriter_l_inst_l_returnflag_o_chars_dvalid,
      l_returnflag_o_chars_last        => PriceSummaryWriter_l_inst_l_returnflag_o_chars_last,
      l_returnflag_o_chars             => PriceSummaryWriter_l_inst_l_returnflag_o_chars,
      l_returnflag_o_chars_count       => PriceSummaryWriter_l_inst_l_returnflag_o_chars_count,
      l_returnflag_o_bus_wreq_valid    => PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_valid,
      l_returnflag_o_bus_wreq_ready    => PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_ready,
      l_returnflag_o_bus_wreq_addr     => PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_addr,
      l_returnflag_o_bus_wreq_len      => PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_len,
      l_returnflag_o_bus_wdat_valid    => PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_valid,
      l_returnflag_o_bus_wdat_ready    => PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_ready,
      l_returnflag_o_bus_wdat_data     => PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_data,
      l_returnflag_o_bus_wdat_strobe   => PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_strobe,
      l_returnflag_o_bus_wdat_last     => PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_last,
      l_returnflag_o_cmd_valid         => PriceSummaryWriter_l_inst_l_returnflag_o_cmd_valid,
      l_returnflag_o_cmd_ready         => PriceSummaryWriter_l_inst_l_returnflag_o_cmd_ready,
      l_returnflag_o_cmd_firstIdx      => PriceSummaryWriter_l_inst_l_returnflag_o_cmd_firstIdx,
      l_returnflag_o_cmd_lastIdx       => PriceSummaryWriter_l_inst_l_returnflag_o_cmd_lastIdx,
      l_returnflag_o_cmd_ctrl          => PriceSummaryWriter_l_inst_l_returnflag_o_cmd_ctrl,
      l_returnflag_o_cmd_tag           => PriceSummaryWriter_l_inst_l_returnflag_o_cmd_tag,
      l_returnflag_o_unl_valid         => PriceSummaryWriter_l_inst_l_returnflag_o_unl_valid,
      l_returnflag_o_unl_ready         => PriceSummaryWriter_l_inst_l_returnflag_o_unl_ready,
      l_returnflag_o_unl_tag           => PriceSummaryWriter_l_inst_l_returnflag_o_unl_tag,
      l_linestatus_o_valid             => PriceSummaryWriter_l_inst_l_linestatus_o_valid,
      l_linestatus_o_ready             => PriceSummaryWriter_l_inst_l_linestatus_o_ready,
      l_linestatus_o_dvalid            => PriceSummaryWriter_l_inst_l_linestatus_o_dvalid,
      l_linestatus_o_last              => PriceSummaryWriter_l_inst_l_linestatus_o_last,
      l_linestatus_o_length            => PriceSummaryWriter_l_inst_l_linestatus_o_length,
      l_linestatus_o_count             => PriceSummaryWriter_l_inst_l_linestatus_o_count,
      l_linestatus_o_chars_valid       => PriceSummaryWriter_l_inst_l_linestatus_o_chars_valid,
      l_linestatus_o_chars_ready       => PriceSummaryWriter_l_inst_l_linestatus_o_chars_ready,
      l_linestatus_o_chars_dvalid      => PriceSummaryWriter_l_inst_l_linestatus_o_chars_dvalid,
      l_linestatus_o_chars_last        => PriceSummaryWriter_l_inst_l_linestatus_o_chars_last,
      l_linestatus_o_chars             => PriceSummaryWriter_l_inst_l_linestatus_o_chars,
      l_linestatus_o_chars_count       => PriceSummaryWriter_l_inst_l_linestatus_o_chars_count,
      l_linestatus_o_bus_wreq_valid    => PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_valid,
      l_linestatus_o_bus_wreq_ready    => PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_ready,
      l_linestatus_o_bus_wreq_addr     => PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_addr,
      l_linestatus_o_bus_wreq_len      => PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_len,
      l_linestatus_o_bus_wdat_valid    => PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_valid,
      l_linestatus_o_bus_wdat_ready    => PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_ready,
      l_linestatus_o_bus_wdat_data     => PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_data,
      l_linestatus_o_bus_wdat_strobe   => PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_strobe,
      l_linestatus_o_bus_wdat_last     => PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_last,
      l_linestatus_o_cmd_valid         => PriceSummaryWriter_l_inst_l_linestatus_o_cmd_valid,
      l_linestatus_o_cmd_ready         => PriceSummaryWriter_l_inst_l_linestatus_o_cmd_ready,
      l_linestatus_o_cmd_firstIdx      => PriceSummaryWriter_l_inst_l_linestatus_o_cmd_firstIdx,
      l_linestatus_o_cmd_lastIdx       => PriceSummaryWriter_l_inst_l_linestatus_o_cmd_lastIdx,
      l_linestatus_o_cmd_ctrl          => PriceSummaryWriter_l_inst_l_linestatus_o_cmd_ctrl,
      l_linestatus_o_cmd_tag           => PriceSummaryWriter_l_inst_l_linestatus_o_cmd_tag,
      l_linestatus_o_unl_valid         => PriceSummaryWriter_l_inst_l_linestatus_o_unl_valid,
      l_linestatus_o_unl_ready         => PriceSummaryWriter_l_inst_l_linestatus_o_unl_ready,
      l_linestatus_o_unl_tag           => PriceSummaryWriter_l_inst_l_linestatus_o_unl_tag,
      l_sum_qty_valid                  => PriceSummaryWriter_l_inst_l_sum_qty_valid,
      l_sum_qty_ready                  => PriceSummaryWriter_l_inst_l_sum_qty_ready,
      l_sum_qty_dvalid                 => PriceSummaryWriter_l_inst_l_sum_qty_dvalid,
      l_sum_qty_last                   => PriceSummaryWriter_l_inst_l_sum_qty_last,
      l_sum_qty                        => PriceSummaryWriter_l_inst_l_sum_qty,
      l_sum_qty_bus_wreq_valid         => PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_valid,
      l_sum_qty_bus_wreq_ready         => PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_ready,
      l_sum_qty_bus_wreq_addr          => PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_addr,
      l_sum_qty_bus_wreq_len           => PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_len,
      l_sum_qty_bus_wdat_valid         => PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_valid,
      l_sum_qty_bus_wdat_ready         => PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_ready,
      l_sum_qty_bus_wdat_data          => PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_data,
      l_sum_qty_bus_wdat_strobe        => PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_strobe,
      l_sum_qty_bus_wdat_last          => PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_last,
      l_sum_qty_cmd_valid              => PriceSummaryWriter_l_inst_l_sum_qty_cmd_valid,
      l_sum_qty_cmd_ready              => PriceSummaryWriter_l_inst_l_sum_qty_cmd_ready,
      l_sum_qty_cmd_firstIdx           => PriceSummaryWriter_l_inst_l_sum_qty_cmd_firstIdx,
      l_sum_qty_cmd_lastIdx            => PriceSummaryWriter_l_inst_l_sum_qty_cmd_lastIdx,
      l_sum_qty_cmd_ctrl               => PriceSummaryWriter_l_inst_l_sum_qty_cmd_ctrl,
      l_sum_qty_cmd_tag                => PriceSummaryWriter_l_inst_l_sum_qty_cmd_tag,
      l_sum_qty_unl_valid              => PriceSummaryWriter_l_inst_l_sum_qty_unl_valid,
      l_sum_qty_unl_ready              => PriceSummaryWriter_l_inst_l_sum_qty_unl_ready,
      l_sum_qty_unl_tag                => PriceSummaryWriter_l_inst_l_sum_qty_unl_tag,
      l_sum_base_price_valid           => PriceSummaryWriter_l_inst_l_sum_base_price_valid,
      l_sum_base_price_ready           => PriceSummaryWriter_l_inst_l_sum_base_price_ready,
      l_sum_base_price_dvalid          => PriceSummaryWriter_l_inst_l_sum_base_price_dvalid,
      l_sum_base_price_last            => PriceSummaryWriter_l_inst_l_sum_base_price_last,
      l_sum_base_price                 => PriceSummaryWriter_l_inst_l_sum_base_price,
      l_sum_base_price_bus_wreq_valid  => PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_valid,
      l_sum_base_price_bus_wreq_ready  => PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_ready,
      l_sum_base_price_bus_wreq_addr   => PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_addr,
      l_sum_base_price_bus_wreq_len    => PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_len,
      l_sum_base_price_bus_wdat_valid  => PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_valid,
      l_sum_base_price_bus_wdat_ready  => PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_ready,
      l_sum_base_price_bus_wdat_data   => PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_data,
      l_sum_base_price_bus_wdat_strobe => PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_strobe,
      l_sum_base_price_bus_wdat_last   => PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_last,
      l_sum_base_price_cmd_valid       => PriceSummaryWriter_l_inst_l_sum_base_price_cmd_valid,
      l_sum_base_price_cmd_ready       => PriceSummaryWriter_l_inst_l_sum_base_price_cmd_ready,
      l_sum_base_price_cmd_firstIdx    => PriceSummaryWriter_l_inst_l_sum_base_price_cmd_firstIdx,
      l_sum_base_price_cmd_lastIdx     => PriceSummaryWriter_l_inst_l_sum_base_price_cmd_lastIdx,
      l_sum_base_price_cmd_ctrl        => PriceSummaryWriter_l_inst_l_sum_base_price_cmd_ctrl,
      l_sum_base_price_cmd_tag         => PriceSummaryWriter_l_inst_l_sum_base_price_cmd_tag,
      l_sum_base_price_unl_valid       => PriceSummaryWriter_l_inst_l_sum_base_price_unl_valid,
      l_sum_base_price_unl_ready       => PriceSummaryWriter_l_inst_l_sum_base_price_unl_ready,
      l_sum_base_price_unl_tag         => PriceSummaryWriter_l_inst_l_sum_base_price_unl_tag,
      l_sum_disc_price_valid           => PriceSummaryWriter_l_inst_l_sum_disc_price_valid,
      l_sum_disc_price_ready           => PriceSummaryWriter_l_inst_l_sum_disc_price_ready,
      l_sum_disc_price_dvalid          => PriceSummaryWriter_l_inst_l_sum_disc_price_dvalid,
      l_sum_disc_price_last            => PriceSummaryWriter_l_inst_l_sum_disc_price_last,
      l_sum_disc_price                 => PriceSummaryWriter_l_inst_l_sum_disc_price,
      l_sum_disc_price_bus_wreq_valid  => PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_valid,
      l_sum_disc_price_bus_wreq_ready  => PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_ready,
      l_sum_disc_price_bus_wreq_addr   => PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_addr,
      l_sum_disc_price_bus_wreq_len    => PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_len,
      l_sum_disc_price_bus_wdat_valid  => PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_valid,
      l_sum_disc_price_bus_wdat_ready  => PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_ready,
      l_sum_disc_price_bus_wdat_data   => PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_data,
      l_sum_disc_price_bus_wdat_strobe => PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_strobe,
      l_sum_disc_price_bus_wdat_last   => PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_last,
      l_sum_disc_price_cmd_valid       => PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_valid,
      l_sum_disc_price_cmd_ready       => PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_ready,
      l_sum_disc_price_cmd_firstIdx    => PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_firstIdx,
      l_sum_disc_price_cmd_lastIdx     => PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_lastIdx,
      l_sum_disc_price_cmd_ctrl        => PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_ctrl,
      l_sum_disc_price_cmd_tag         => PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_tag,
      l_sum_disc_price_unl_valid       => PriceSummaryWriter_l_inst_l_sum_disc_price_unl_valid,
      l_sum_disc_price_unl_ready       => PriceSummaryWriter_l_inst_l_sum_disc_price_unl_ready,
      l_sum_disc_price_unl_tag         => PriceSummaryWriter_l_inst_l_sum_disc_price_unl_tag,
      l_sum_charge_valid               => PriceSummaryWriter_l_inst_l_sum_charge_valid,
      l_sum_charge_ready               => PriceSummaryWriter_l_inst_l_sum_charge_ready,
      l_sum_charge_dvalid              => PriceSummaryWriter_l_inst_l_sum_charge_dvalid,
      l_sum_charge_last                => PriceSummaryWriter_l_inst_l_sum_charge_last,
      l_sum_charge                     => PriceSummaryWriter_l_inst_l_sum_charge,
      l_sum_charge_bus_wreq_valid      => PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_valid,
      l_sum_charge_bus_wreq_ready      => PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_ready,
      l_sum_charge_bus_wreq_addr       => PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_addr,
      l_sum_charge_bus_wreq_len        => PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_len,
      l_sum_charge_bus_wdat_valid      => PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_valid,
      l_sum_charge_bus_wdat_ready      => PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_ready,
      l_sum_charge_bus_wdat_data       => PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_data,
      l_sum_charge_bus_wdat_strobe     => PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_strobe,
      l_sum_charge_bus_wdat_last       => PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_last,
      l_sum_charge_cmd_valid           => PriceSummaryWriter_l_inst_l_sum_charge_cmd_valid,
      l_sum_charge_cmd_ready           => PriceSummaryWriter_l_inst_l_sum_charge_cmd_ready,
      l_sum_charge_cmd_firstIdx        => PriceSummaryWriter_l_inst_l_sum_charge_cmd_firstIdx,
      l_sum_charge_cmd_lastIdx         => PriceSummaryWriter_l_inst_l_sum_charge_cmd_lastIdx,
      l_sum_charge_cmd_ctrl            => PriceSummaryWriter_l_inst_l_sum_charge_cmd_ctrl,
      l_sum_charge_cmd_tag             => PriceSummaryWriter_l_inst_l_sum_charge_cmd_tag,
      l_sum_charge_unl_valid           => PriceSummaryWriter_l_inst_l_sum_charge_unl_valid,
      l_sum_charge_unl_ready           => PriceSummaryWriter_l_inst_l_sum_charge_unl_ready,
      l_sum_charge_unl_tag             => PriceSummaryWriter_l_inst_l_sum_charge_unl_tag,
      l_avg_qty_valid                  => PriceSummaryWriter_l_inst_l_avg_qty_valid,
      l_avg_qty_ready                  => PriceSummaryWriter_l_inst_l_avg_qty_ready,
      l_avg_qty_dvalid                 => PriceSummaryWriter_l_inst_l_avg_qty_dvalid,
      l_avg_qty_last                   => PriceSummaryWriter_l_inst_l_avg_qty_last,
      l_avg_qty                        => PriceSummaryWriter_l_inst_l_avg_qty,
      l_avg_qty_bus_wreq_valid         => PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_valid,
      l_avg_qty_bus_wreq_ready         => PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_ready,
      l_avg_qty_bus_wreq_addr          => PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_addr,
      l_avg_qty_bus_wreq_len           => PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_len,
      l_avg_qty_bus_wdat_valid         => PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_valid,
      l_avg_qty_bus_wdat_ready         => PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_ready,
      l_avg_qty_bus_wdat_data          => PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_data,
      l_avg_qty_bus_wdat_strobe        => PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_strobe,
      l_avg_qty_bus_wdat_last          => PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_last,
      l_avg_qty_cmd_valid              => PriceSummaryWriter_l_inst_l_avg_qty_cmd_valid,
      l_avg_qty_cmd_ready              => PriceSummaryWriter_l_inst_l_avg_qty_cmd_ready,
      l_avg_qty_cmd_firstIdx           => PriceSummaryWriter_l_inst_l_avg_qty_cmd_firstIdx,
      l_avg_qty_cmd_lastIdx            => PriceSummaryWriter_l_inst_l_avg_qty_cmd_lastIdx,
      l_avg_qty_cmd_ctrl               => PriceSummaryWriter_l_inst_l_avg_qty_cmd_ctrl,
      l_avg_qty_cmd_tag                => PriceSummaryWriter_l_inst_l_avg_qty_cmd_tag,
      l_avg_qty_unl_valid              => PriceSummaryWriter_l_inst_l_avg_qty_unl_valid,
      l_avg_qty_unl_ready              => PriceSummaryWriter_l_inst_l_avg_qty_unl_ready,
      l_avg_qty_unl_tag                => PriceSummaryWriter_l_inst_l_avg_qty_unl_tag,
      l_avg_price_valid                => PriceSummaryWriter_l_inst_l_avg_price_valid,
      l_avg_price_ready                => PriceSummaryWriter_l_inst_l_avg_price_ready,
      l_avg_price_dvalid               => PriceSummaryWriter_l_inst_l_avg_price_dvalid,
      l_avg_price_last                 => PriceSummaryWriter_l_inst_l_avg_price_last,
      l_avg_price                      => PriceSummaryWriter_l_inst_l_avg_price,
      l_avg_price_bus_wreq_valid       => PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_valid,
      l_avg_price_bus_wreq_ready       => PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_ready,
      l_avg_price_bus_wreq_addr        => PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_addr,
      l_avg_price_bus_wreq_len         => PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_len,
      l_avg_price_bus_wdat_valid       => PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_valid,
      l_avg_price_bus_wdat_ready       => PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_ready,
      l_avg_price_bus_wdat_data        => PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_data,
      l_avg_price_bus_wdat_strobe      => PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_strobe,
      l_avg_price_bus_wdat_last        => PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_last,
      l_avg_price_cmd_valid            => PriceSummaryWriter_l_inst_l_avg_price_cmd_valid,
      l_avg_price_cmd_ready            => PriceSummaryWriter_l_inst_l_avg_price_cmd_ready,
      l_avg_price_cmd_firstIdx         => PriceSummaryWriter_l_inst_l_avg_price_cmd_firstIdx,
      l_avg_price_cmd_lastIdx          => PriceSummaryWriter_l_inst_l_avg_price_cmd_lastIdx,
      l_avg_price_cmd_ctrl             => PriceSummaryWriter_l_inst_l_avg_price_cmd_ctrl,
      l_avg_price_cmd_tag              => PriceSummaryWriter_l_inst_l_avg_price_cmd_tag,
      l_avg_price_unl_valid            => PriceSummaryWriter_l_inst_l_avg_price_unl_valid,
      l_avg_price_unl_ready            => PriceSummaryWriter_l_inst_l_avg_price_unl_ready,
      l_avg_price_unl_tag              => PriceSummaryWriter_l_inst_l_avg_price_unl_tag,
      l_avg_disc_valid                 => PriceSummaryWriter_l_inst_l_avg_disc_valid,
      l_avg_disc_ready                 => PriceSummaryWriter_l_inst_l_avg_disc_ready,
      l_avg_disc_dvalid                => PriceSummaryWriter_l_inst_l_avg_disc_dvalid,
      l_avg_disc_last                  => PriceSummaryWriter_l_inst_l_avg_disc_last,
      l_avg_disc                       => PriceSummaryWriter_l_inst_l_avg_disc,
      l_avg_disc_bus_wreq_valid        => PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_valid,
      l_avg_disc_bus_wreq_ready        => PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_ready,
      l_avg_disc_bus_wreq_addr         => PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_addr,
      l_avg_disc_bus_wreq_len          => PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_len,
      l_avg_disc_bus_wdat_valid        => PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_valid,
      l_avg_disc_bus_wdat_ready        => PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_ready,
      l_avg_disc_bus_wdat_data         => PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_data,
      l_avg_disc_bus_wdat_strobe       => PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_strobe,
      l_avg_disc_bus_wdat_last         => PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_last,
      l_avg_disc_cmd_valid             => PriceSummaryWriter_l_inst_l_avg_disc_cmd_valid,
      l_avg_disc_cmd_ready             => PriceSummaryWriter_l_inst_l_avg_disc_cmd_ready,
      l_avg_disc_cmd_firstIdx          => PriceSummaryWriter_l_inst_l_avg_disc_cmd_firstIdx,
      l_avg_disc_cmd_lastIdx           => PriceSummaryWriter_l_inst_l_avg_disc_cmd_lastIdx,
      l_avg_disc_cmd_ctrl              => PriceSummaryWriter_l_inst_l_avg_disc_cmd_ctrl,
      l_avg_disc_cmd_tag               => PriceSummaryWriter_l_inst_l_avg_disc_cmd_tag,
      l_avg_disc_unl_valid             => PriceSummaryWriter_l_inst_l_avg_disc_unl_valid,
      l_avg_disc_unl_ready             => PriceSummaryWriter_l_inst_l_avg_disc_unl_ready,
      l_avg_disc_unl_tag               => PriceSummaryWriter_l_inst_l_avg_disc_unl_tag,
      l_count_order_valid              => PriceSummaryWriter_l_inst_l_count_order_valid,
      l_count_order_ready              => PriceSummaryWriter_l_inst_l_count_order_ready,
      l_count_order_dvalid             => PriceSummaryWriter_l_inst_l_count_order_dvalid,
      l_count_order_last               => PriceSummaryWriter_l_inst_l_count_order_last,
      l_count_order                    => PriceSummaryWriter_l_inst_l_count_order,
      l_count_order_bus_wreq_valid     => PriceSummaryWriter_l_inst_l_count_order_bus_wreq_valid,
      l_count_order_bus_wreq_ready     => PriceSummaryWriter_l_inst_l_count_order_bus_wreq_ready,
      l_count_order_bus_wreq_addr      => PriceSummaryWriter_l_inst_l_count_order_bus_wreq_addr,
      l_count_order_bus_wreq_len       => PriceSummaryWriter_l_inst_l_count_order_bus_wreq_len,
      l_count_order_bus_wdat_valid     => PriceSummaryWriter_l_inst_l_count_order_bus_wdat_valid,
      l_count_order_bus_wdat_ready     => PriceSummaryWriter_l_inst_l_count_order_bus_wdat_ready,
      l_count_order_bus_wdat_data      => PriceSummaryWriter_l_inst_l_count_order_bus_wdat_data,
      l_count_order_bus_wdat_strobe    => PriceSummaryWriter_l_inst_l_count_order_bus_wdat_strobe,
      l_count_order_bus_wdat_last      => PriceSummaryWriter_l_inst_l_count_order_bus_wdat_last,
      l_count_order_cmd_valid          => PriceSummaryWriter_l_inst_l_count_order_cmd_valid,
      l_count_order_cmd_ready          => PriceSummaryWriter_l_inst_l_count_order_cmd_ready,
      l_count_order_cmd_firstIdx       => PriceSummaryWriter_l_inst_l_count_order_cmd_firstIdx,
      l_count_order_cmd_lastIdx        => PriceSummaryWriter_l_inst_l_count_order_cmd_lastIdx,
      l_count_order_cmd_ctrl           => PriceSummaryWriter_l_inst_l_count_order_cmd_ctrl,
      l_count_order_cmd_tag            => PriceSummaryWriter_l_inst_l_count_order_cmd_tag,
      l_count_order_unl_valid          => PriceSummaryWriter_l_inst_l_count_order_unl_valid,
      l_count_order_unl_ready          => PriceSummaryWriter_l_inst_l_count_order_unl_ready,
      l_count_order_unl_tag            => PriceSummaryWriter_l_inst_l_count_order_unl_tag
    );

  WRAW64DW512LW8BS1BM16_inst : BusWriteArbiterVec
    generic map (
      BUS_ADDR_WIDTH  => BUS_ADDR_WIDTH,
      BUS_DATA_WIDTH  => BUS_DATA_WIDTH,
      BUS_LEN_WIDTH   => BUS_LEN_WIDTH,
      NUM_SLAVE_PORTS => 10,
      ARB_METHOD      => "RR-STICKY",
      MAX_OUTSTANDING => 4,
      RAM_CONFIG      => "",
      SLV_REQ_SLICES  => true,
      MST_REQ_SLICE   => true,
      MST_DAT_SLICE   => true,
      SLV_DAT_SLICES  => true
    )
    port map (
      bcd_clk         => bcd_clk,
      bcd_reset       => bcd_reset,
      mst_wreq_valid  => WRAW64DW512LW8BS1BM16_inst_mst_wreq_valid,
      mst_wreq_ready  => WRAW64DW512LW8BS1BM16_inst_mst_wreq_ready,
      mst_wreq_addr   => WRAW64DW512LW8BS1BM16_inst_mst_wreq_addr,
      mst_wreq_len    => WRAW64DW512LW8BS1BM16_inst_mst_wreq_len,
      mst_wdat_valid  => WRAW64DW512LW8BS1BM16_inst_mst_wdat_valid,
      mst_wdat_ready  => WRAW64DW512LW8BS1BM16_inst_mst_wdat_ready,
      mst_wdat_data   => WRAW64DW512LW8BS1BM16_inst_mst_wdat_data,
      mst_wdat_strobe => WRAW64DW512LW8BS1BM16_inst_mst_wdat_strobe,
      mst_wdat_last   => WRAW64DW512LW8BS1BM16_inst_mst_wdat_last,
      bsv_wreq_valid  => WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid,
      bsv_wreq_ready  => WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready,
      bsv_wreq_len    => WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len,
      bsv_wreq_addr   => WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr,
      bsv_wdat_valid  => WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid,
      bsv_wdat_strobe => WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe,
      bsv_wdat_ready  => WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready,
      bsv_wdat_last   => WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last,
      bsv_wdat_data   => WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data
    );

  wr_mst_wreq_valid                         <= WRAW64DW512LW8BS1BM16_inst_mst_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_mst_wreq_ready <= wr_mst_wreq_ready;
  wr_mst_wreq_addr                          <= WRAW64DW512LW8BS1BM16_inst_mst_wreq_addr;
  wr_mst_wreq_len                           <= WRAW64DW512LW8BS1BM16_inst_mst_wreq_len;
  wr_mst_wdat_valid                         <= WRAW64DW512LW8BS1BM16_inst_mst_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_mst_wdat_ready <= wr_mst_wdat_ready;
  wr_mst_wdat_data                          <= WRAW64DW512LW8BS1BM16_inst_mst_wdat_data;
  wr_mst_wdat_strobe                        <= WRAW64DW512LW8BS1BM16_inst_mst_wdat_strobe;
  wr_mst_wdat_last                          <= WRAW64DW512LW8BS1BM16_inst_mst_wdat_last;

  PriceSummaryWriter_Nucleus_inst_mmio_awvalid               <= mmio_awvalid;
  mmio_awready                                               <= PriceSummaryWriter_Nucleus_inst_mmio_awready;
  PriceSummaryWriter_Nucleus_inst_mmio_awaddr                <= mmio_awaddr;
  PriceSummaryWriter_Nucleus_inst_mmio_wvalid                <= mmio_wvalid;
  mmio_wready                                                <= PriceSummaryWriter_Nucleus_inst_mmio_wready;
  PriceSummaryWriter_Nucleus_inst_mmio_wdata                 <= mmio_wdata;
  PriceSummaryWriter_Nucleus_inst_mmio_wstrb                 <= mmio_wstrb;
  mmio_bvalid                                                <= PriceSummaryWriter_Nucleus_inst_mmio_bvalid;
  PriceSummaryWriter_Nucleus_inst_mmio_bready                <= mmio_bready;
  mmio_bresp                                                 <= PriceSummaryWriter_Nucleus_inst_mmio_bresp;
  PriceSummaryWriter_Nucleus_inst_mmio_arvalid               <= mmio_arvalid;
  mmio_arready                                               <= PriceSummaryWriter_Nucleus_inst_mmio_arready;
  PriceSummaryWriter_Nucleus_inst_mmio_araddr                <= mmio_araddr;
  mmio_rvalid                                                <= PriceSummaryWriter_Nucleus_inst_mmio_rvalid;
  PriceSummaryWriter_Nucleus_inst_mmio_rready                <= mmio_rready;
  mmio_rdata                                                 <= PriceSummaryWriter_Nucleus_inst_mmio_rdata;
  mmio_rresp                                                 <= PriceSummaryWriter_Nucleus_inst_mmio_rresp;

  PriceSummaryWriter_Nucleus_inst_l_returnflag_o_unl_valid   <= PriceSummaryWriter_l_inst_l_returnflag_o_unl_valid;
  PriceSummaryWriter_l_inst_l_returnflag_o_unl_ready         <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_unl_ready;
  PriceSummaryWriter_Nucleus_inst_l_returnflag_o_unl_tag     <= PriceSummaryWriter_l_inst_l_returnflag_o_unl_tag;

  PriceSummaryWriter_Nucleus_inst_l_linestatus_o_unl_valid   <= PriceSummaryWriter_l_inst_l_linestatus_o_unl_valid;
  PriceSummaryWriter_l_inst_l_linestatus_o_unl_ready         <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_unl_ready;
  PriceSummaryWriter_Nucleus_inst_l_linestatus_o_unl_tag     <= PriceSummaryWriter_l_inst_l_linestatus_o_unl_tag;

  PriceSummaryWriter_Nucleus_inst_l_sum_qty_unl_valid        <= PriceSummaryWriter_l_inst_l_sum_qty_unl_valid;
  PriceSummaryWriter_l_inst_l_sum_qty_unl_ready              <= PriceSummaryWriter_Nucleus_inst_l_sum_qty_unl_ready;
  PriceSummaryWriter_Nucleus_inst_l_sum_qty_unl_tag          <= PriceSummaryWriter_l_inst_l_sum_qty_unl_tag;

  PriceSummaryWriter_Nucleus_inst_l_sum_base_price_unl_valid <= PriceSummaryWriter_l_inst_l_sum_base_price_unl_valid;
  PriceSummaryWriter_l_inst_l_sum_base_price_unl_ready       <= PriceSummaryWriter_Nucleus_inst_l_sum_base_price_unl_ready;
  PriceSummaryWriter_Nucleus_inst_l_sum_base_price_unl_tag   <= PriceSummaryWriter_l_inst_l_sum_base_price_unl_tag;

  PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_unl_valid <= PriceSummaryWriter_l_inst_l_sum_disc_price_unl_valid;
  PriceSummaryWriter_l_inst_l_sum_disc_price_unl_ready       <= PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_unl_ready;
  PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_unl_tag   <= PriceSummaryWriter_l_inst_l_sum_disc_price_unl_tag;

  PriceSummaryWriter_Nucleus_inst_l_sum_charge_unl_valid     <= PriceSummaryWriter_l_inst_l_sum_charge_unl_valid;
  PriceSummaryWriter_l_inst_l_sum_charge_unl_ready           <= PriceSummaryWriter_Nucleus_inst_l_sum_charge_unl_ready;
  PriceSummaryWriter_Nucleus_inst_l_sum_charge_unl_tag       <= PriceSummaryWriter_l_inst_l_sum_charge_unl_tag;

  PriceSummaryWriter_Nucleus_inst_l_avg_qty_unl_valid        <= PriceSummaryWriter_l_inst_l_avg_qty_unl_valid;
  PriceSummaryWriter_l_inst_l_avg_qty_unl_ready              <= PriceSummaryWriter_Nucleus_inst_l_avg_qty_unl_ready;
  PriceSummaryWriter_Nucleus_inst_l_avg_qty_unl_tag          <= PriceSummaryWriter_l_inst_l_avg_qty_unl_tag;

  PriceSummaryWriter_Nucleus_inst_l_avg_price_unl_valid      <= PriceSummaryWriter_l_inst_l_avg_price_unl_valid;
  PriceSummaryWriter_l_inst_l_avg_price_unl_ready            <= PriceSummaryWriter_Nucleus_inst_l_avg_price_unl_ready;
  PriceSummaryWriter_Nucleus_inst_l_avg_price_unl_tag        <= PriceSummaryWriter_l_inst_l_avg_price_unl_tag;

  PriceSummaryWriter_Nucleus_inst_l_avg_disc_unl_valid       <= PriceSummaryWriter_l_inst_l_avg_disc_unl_valid;
  PriceSummaryWriter_l_inst_l_avg_disc_unl_ready             <= PriceSummaryWriter_Nucleus_inst_l_avg_disc_unl_ready;
  PriceSummaryWriter_Nucleus_inst_l_avg_disc_unl_tag         <= PriceSummaryWriter_l_inst_l_avg_disc_unl_tag;

  PriceSummaryWriter_Nucleus_inst_l_count_order_unl_valid    <= PriceSummaryWriter_l_inst_l_count_order_unl_valid;
  PriceSummaryWriter_l_inst_l_count_order_unl_ready          <= PriceSummaryWriter_Nucleus_inst_l_count_order_unl_ready;
  PriceSummaryWriter_Nucleus_inst_l_count_order_unl_tag      <= PriceSummaryWriter_l_inst_l_count_order_unl_tag;

  PriceSummaryWriter_l_inst_l_returnflag_o_valid             <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_valid;
  PriceSummaryWriter_Nucleus_inst_l_returnflag_o_ready       <= PriceSummaryWriter_l_inst_l_returnflag_o_ready;
  PriceSummaryWriter_l_inst_l_returnflag_o_dvalid            <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_dvalid;
  PriceSummaryWriter_l_inst_l_returnflag_o_last              <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_last;
  PriceSummaryWriter_l_inst_l_returnflag_o_length            <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_length;
  PriceSummaryWriter_l_inst_l_returnflag_o_count             <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_count;
  PriceSummaryWriter_l_inst_l_returnflag_o_chars_valid       <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_valid;
  PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_ready <= PriceSummaryWriter_l_inst_l_returnflag_o_chars_ready;
  PriceSummaryWriter_l_inst_l_returnflag_o_chars_dvalid      <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_dvalid;
  PriceSummaryWriter_l_inst_l_returnflag_o_chars_last        <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_last;
  PriceSummaryWriter_l_inst_l_returnflag_o_chars             <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars;
  PriceSummaryWriter_l_inst_l_returnflag_o_chars_count       <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_chars_count;

  PriceSummaryWriter_l_inst_l_returnflag_o_cmd_valid         <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_valid;
  PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_ready   <= PriceSummaryWriter_l_inst_l_returnflag_o_cmd_ready;
  PriceSummaryWriter_l_inst_l_returnflag_o_cmd_firstIdx      <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_firstIdx;
  PriceSummaryWriter_l_inst_l_returnflag_o_cmd_lastIdx       <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_lastIdx;
  PriceSummaryWriter_l_inst_l_returnflag_o_cmd_ctrl          <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_ctrl;
  PriceSummaryWriter_l_inst_l_returnflag_o_cmd_tag           <= PriceSummaryWriter_Nucleus_inst_l_returnflag_o_cmd_tag;

  PriceSummaryWriter_l_inst_l_linestatus_o_valid             <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_valid;
  PriceSummaryWriter_Nucleus_inst_l_linestatus_o_ready       <= PriceSummaryWriter_l_inst_l_linestatus_o_ready;
  PriceSummaryWriter_l_inst_l_linestatus_o_dvalid            <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_dvalid;
  PriceSummaryWriter_l_inst_l_linestatus_o_last              <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_last;
  PriceSummaryWriter_l_inst_l_linestatus_o_length            <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_length;
  PriceSummaryWriter_l_inst_l_linestatus_o_count             <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_count;
  PriceSummaryWriter_l_inst_l_linestatus_o_chars_valid       <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_valid;
  PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_ready <= PriceSummaryWriter_l_inst_l_linestatus_o_chars_ready;
  PriceSummaryWriter_l_inst_l_linestatus_o_chars_dvalid      <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_dvalid;
  PriceSummaryWriter_l_inst_l_linestatus_o_chars_last        <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_last;
  PriceSummaryWriter_l_inst_l_linestatus_o_chars             <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars;
  PriceSummaryWriter_l_inst_l_linestatus_o_chars_count       <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_chars_count;

  PriceSummaryWriter_l_inst_l_linestatus_o_cmd_valid         <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_valid;
  PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_ready   <= PriceSummaryWriter_l_inst_l_linestatus_o_cmd_ready;
  PriceSummaryWriter_l_inst_l_linestatus_o_cmd_firstIdx      <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_firstIdx;
  PriceSummaryWriter_l_inst_l_linestatus_o_cmd_lastIdx       <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_lastIdx;
  PriceSummaryWriter_l_inst_l_linestatus_o_cmd_ctrl          <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_ctrl;
  PriceSummaryWriter_l_inst_l_linestatus_o_cmd_tag           <= PriceSummaryWriter_Nucleus_inst_l_linestatus_o_cmd_tag;

  PriceSummaryWriter_l_inst_l_sum_qty_valid                  <= PriceSummaryWriter_Nucleus_inst_l_sum_qty_valid;
  PriceSummaryWriter_Nucleus_inst_l_sum_qty_ready            <= PriceSummaryWriter_l_inst_l_sum_qty_ready;
  PriceSummaryWriter_l_inst_l_sum_qty_dvalid                 <= PriceSummaryWriter_Nucleus_inst_l_sum_qty_dvalid;
  PriceSummaryWriter_l_inst_l_sum_qty_last                   <= PriceSummaryWriter_Nucleus_inst_l_sum_qty_last;
  PriceSummaryWriter_l_inst_l_sum_qty                        <= PriceSummaryWriter_Nucleus_inst_l_sum_qty;

  PriceSummaryWriter_l_inst_l_sum_qty_cmd_valid              <= PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_valid;
  PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_ready        <= PriceSummaryWriter_l_inst_l_sum_qty_cmd_ready;
  PriceSummaryWriter_l_inst_l_sum_qty_cmd_firstIdx           <= PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_firstIdx;
  PriceSummaryWriter_l_inst_l_sum_qty_cmd_lastIdx            <= PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_lastIdx;
  PriceSummaryWriter_l_inst_l_sum_qty_cmd_ctrl               <= PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_ctrl;
  PriceSummaryWriter_l_inst_l_sum_qty_cmd_tag                <= PriceSummaryWriter_Nucleus_inst_l_sum_qty_cmd_tag;

  PriceSummaryWriter_l_inst_l_sum_base_price_valid           <= PriceSummaryWriter_Nucleus_inst_l_sum_base_price_valid;
  PriceSummaryWriter_Nucleus_inst_l_sum_base_price_ready     <= PriceSummaryWriter_l_inst_l_sum_base_price_ready;
  PriceSummaryWriter_l_inst_l_sum_base_price_dvalid          <= PriceSummaryWriter_Nucleus_inst_l_sum_base_price_dvalid;
  PriceSummaryWriter_l_inst_l_sum_base_price_last            <= PriceSummaryWriter_Nucleus_inst_l_sum_base_price_last;
  PriceSummaryWriter_l_inst_l_sum_base_price                 <= PriceSummaryWriter_Nucleus_inst_l_sum_base_price;

  PriceSummaryWriter_l_inst_l_sum_base_price_cmd_valid       <= PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_valid;
  PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_ready <= PriceSummaryWriter_l_inst_l_sum_base_price_cmd_ready;
  PriceSummaryWriter_l_inst_l_sum_base_price_cmd_firstIdx    <= PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_firstIdx;
  PriceSummaryWriter_l_inst_l_sum_base_price_cmd_lastIdx     <= PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_lastIdx;
  PriceSummaryWriter_l_inst_l_sum_base_price_cmd_ctrl        <= PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_ctrl;
  PriceSummaryWriter_l_inst_l_sum_base_price_cmd_tag         <= PriceSummaryWriter_Nucleus_inst_l_sum_base_price_cmd_tag;

  PriceSummaryWriter_l_inst_l_sum_disc_price_valid           <= PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_valid;
  PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_ready     <= PriceSummaryWriter_l_inst_l_sum_disc_price_ready;
  PriceSummaryWriter_l_inst_l_sum_disc_price_dvalid          <= PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_dvalid;
  PriceSummaryWriter_l_inst_l_sum_disc_price_last            <= PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_last;
  PriceSummaryWriter_l_inst_l_sum_disc_price                 <= PriceSummaryWriter_Nucleus_inst_l_sum_disc_price;

  PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_valid       <= PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_valid;
  PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_ready <= PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_ready;
  PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_firstIdx    <= PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_firstIdx;
  PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_lastIdx     <= PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_lastIdx;
  PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_ctrl        <= PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_ctrl;
  PriceSummaryWriter_l_inst_l_sum_disc_price_cmd_tag         <= PriceSummaryWriter_Nucleus_inst_l_sum_disc_price_cmd_tag;

  PriceSummaryWriter_l_inst_l_sum_charge_valid               <= PriceSummaryWriter_Nucleus_inst_l_sum_charge_valid;
  PriceSummaryWriter_Nucleus_inst_l_sum_charge_ready         <= PriceSummaryWriter_l_inst_l_sum_charge_ready;
  PriceSummaryWriter_l_inst_l_sum_charge_dvalid              <= PriceSummaryWriter_Nucleus_inst_l_sum_charge_dvalid;
  PriceSummaryWriter_l_inst_l_sum_charge_last                <= PriceSummaryWriter_Nucleus_inst_l_sum_charge_last;
  PriceSummaryWriter_l_inst_l_sum_charge                     <= PriceSummaryWriter_Nucleus_inst_l_sum_charge;

  PriceSummaryWriter_l_inst_l_sum_charge_cmd_valid           <= PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_valid;
  PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_ready     <= PriceSummaryWriter_l_inst_l_sum_charge_cmd_ready;
  PriceSummaryWriter_l_inst_l_sum_charge_cmd_firstIdx        <= PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_firstIdx;
  PriceSummaryWriter_l_inst_l_sum_charge_cmd_lastIdx         <= PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_lastIdx;
  PriceSummaryWriter_l_inst_l_sum_charge_cmd_ctrl            <= PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_ctrl;
  PriceSummaryWriter_l_inst_l_sum_charge_cmd_tag             <= PriceSummaryWriter_Nucleus_inst_l_sum_charge_cmd_tag;

  PriceSummaryWriter_l_inst_l_avg_qty_valid                  <= PriceSummaryWriter_Nucleus_inst_l_avg_qty_valid;
  PriceSummaryWriter_Nucleus_inst_l_avg_qty_ready            <= PriceSummaryWriter_l_inst_l_avg_qty_ready;
  PriceSummaryWriter_l_inst_l_avg_qty_dvalid                 <= PriceSummaryWriter_Nucleus_inst_l_avg_qty_dvalid;
  PriceSummaryWriter_l_inst_l_avg_qty_last                   <= PriceSummaryWriter_Nucleus_inst_l_avg_qty_last;
  PriceSummaryWriter_l_inst_l_avg_qty                        <= PriceSummaryWriter_Nucleus_inst_l_avg_qty;

  PriceSummaryWriter_l_inst_l_avg_qty_cmd_valid              <= PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_valid;
  PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_ready        <= PriceSummaryWriter_l_inst_l_avg_qty_cmd_ready;
  PriceSummaryWriter_l_inst_l_avg_qty_cmd_firstIdx           <= PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_firstIdx;
  PriceSummaryWriter_l_inst_l_avg_qty_cmd_lastIdx            <= PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_lastIdx;
  PriceSummaryWriter_l_inst_l_avg_qty_cmd_ctrl               <= PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_ctrl;
  PriceSummaryWriter_l_inst_l_avg_qty_cmd_tag                <= PriceSummaryWriter_Nucleus_inst_l_avg_qty_cmd_tag;

  PriceSummaryWriter_l_inst_l_avg_price_valid                <= PriceSummaryWriter_Nucleus_inst_l_avg_price_valid;
  PriceSummaryWriter_Nucleus_inst_l_avg_price_ready          <= PriceSummaryWriter_l_inst_l_avg_price_ready;
  PriceSummaryWriter_l_inst_l_avg_price_dvalid               <= PriceSummaryWriter_Nucleus_inst_l_avg_price_dvalid;
  PriceSummaryWriter_l_inst_l_avg_price_last                 <= PriceSummaryWriter_Nucleus_inst_l_avg_price_last;
  PriceSummaryWriter_l_inst_l_avg_price                      <= PriceSummaryWriter_Nucleus_inst_l_avg_price;

  PriceSummaryWriter_l_inst_l_avg_price_cmd_valid            <= PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_valid;
  PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_ready      <= PriceSummaryWriter_l_inst_l_avg_price_cmd_ready;
  PriceSummaryWriter_l_inst_l_avg_price_cmd_firstIdx         <= PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_firstIdx;
  PriceSummaryWriter_l_inst_l_avg_price_cmd_lastIdx          <= PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_lastIdx;
  PriceSummaryWriter_l_inst_l_avg_price_cmd_ctrl             <= PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_ctrl;
  PriceSummaryWriter_l_inst_l_avg_price_cmd_tag              <= PriceSummaryWriter_Nucleus_inst_l_avg_price_cmd_tag;

  PriceSummaryWriter_l_inst_l_avg_disc_valid                 <= PriceSummaryWriter_Nucleus_inst_l_avg_disc_valid;
  PriceSummaryWriter_Nucleus_inst_l_avg_disc_ready           <= PriceSummaryWriter_l_inst_l_avg_disc_ready;
  PriceSummaryWriter_l_inst_l_avg_disc_dvalid                <= PriceSummaryWriter_Nucleus_inst_l_avg_disc_dvalid;
  PriceSummaryWriter_l_inst_l_avg_disc_last                  <= PriceSummaryWriter_Nucleus_inst_l_avg_disc_last;
  PriceSummaryWriter_l_inst_l_avg_disc                       <= PriceSummaryWriter_Nucleus_inst_l_avg_disc;

  PriceSummaryWriter_l_inst_l_avg_disc_cmd_valid             <= PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_valid;
  PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_ready       <= PriceSummaryWriter_l_inst_l_avg_disc_cmd_ready;
  PriceSummaryWriter_l_inst_l_avg_disc_cmd_firstIdx          <= PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_firstIdx;
  PriceSummaryWriter_l_inst_l_avg_disc_cmd_lastIdx           <= PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_lastIdx;
  PriceSummaryWriter_l_inst_l_avg_disc_cmd_ctrl              <= PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_ctrl;
  PriceSummaryWriter_l_inst_l_avg_disc_cmd_tag               <= PriceSummaryWriter_Nucleus_inst_l_avg_disc_cmd_tag;

  PriceSummaryWriter_l_inst_l_count_order_valid              <= PriceSummaryWriter_Nucleus_inst_l_count_order_valid;
  PriceSummaryWriter_Nucleus_inst_l_count_order_ready        <= PriceSummaryWriter_l_inst_l_count_order_ready;
  PriceSummaryWriter_l_inst_l_count_order_dvalid             <= PriceSummaryWriter_Nucleus_inst_l_count_order_dvalid;
  PriceSummaryWriter_l_inst_l_count_order_last               <= PriceSummaryWriter_Nucleus_inst_l_count_order_last;
  PriceSummaryWriter_l_inst_l_count_order                    <= PriceSummaryWriter_Nucleus_inst_l_count_order;

  PriceSummaryWriter_l_inst_l_count_order_cmd_valid          <= PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_valid;
  PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_ready    <= PriceSummaryWriter_l_inst_l_count_order_cmd_ready;
  PriceSummaryWriter_l_inst_l_count_order_cmd_firstIdx       <= PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_firstIdx;
  PriceSummaryWriter_l_inst_l_count_order_cmd_lastIdx        <= PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_lastIdx;
  PriceSummaryWriter_l_inst_l_count_order_cmd_ctrl           <= PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_ctrl;
  PriceSummaryWriter_l_inst_l_count_order_cmd_tag            <= PriceSummaryWriter_Nucleus_inst_l_count_order_cmd_tag;

  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid(0)                                                                <= PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid(1)                                                                <= PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid(2)                                                                <= PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid(3)                                                                <= PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid(4)                                                                <= PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid(5)                                                                <= PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid(6)                                                                <= PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid(7)                                                                <= PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid(8)                                                                <= PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_valid(9)                                                                <= PriceSummaryWriter_l_inst_l_count_order_bus_wreq_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len(BUS_LEN_WIDTH-1 downto 0)                                           <= PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_len;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len(BUS_LEN_WIDTH+BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH)                 <= PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_len;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len(BUS_LEN_WIDTH*2+BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH*2)             <= PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_len;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len(BUS_LEN_WIDTH*3+BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH*3)             <= PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_len;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len(BUS_LEN_WIDTH*4+BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH*4)             <= PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_len;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len(BUS_LEN_WIDTH*5+BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH*5)             <= PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_len;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len(BUS_LEN_WIDTH*6+BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH*6)             <= PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_len;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len(BUS_LEN_WIDTH*7+BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH*7)             <= PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_len;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len(BUS_LEN_WIDTH*8+BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH*8)             <= PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_len;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_len(BUS_LEN_WIDTH*9+BUS_LEN_WIDTH-1 downto BUS_LEN_WIDTH*9)             <= PriceSummaryWriter_l_inst_l_count_order_bus_wreq_len;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr(BUS_ADDR_WIDTH-1 downto 0)                                         <= PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_addr;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr(BUS_ADDR_WIDTH+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH)             <= PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_addr;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr(BUS_ADDR_WIDTH*2+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH*2)         <= PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_addr;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr(BUS_ADDR_WIDTH*3+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH*3)         <= PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_addr;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr(BUS_ADDR_WIDTH*4+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH*4)         <= PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_addr;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr(BUS_ADDR_WIDTH*5+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH*5)         <= PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_addr;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr(BUS_ADDR_WIDTH*6+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH*6)         <= PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_addr;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr(BUS_ADDR_WIDTH*7+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH*7)         <= PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_addr;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr(BUS_ADDR_WIDTH*8+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH*8)         <= PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_addr;
  WRAW64DW512LW8BS1BM16_inst_bsv_wreq_addr(BUS_ADDR_WIDTH*9+BUS_ADDR_WIDTH-1 downto BUS_ADDR_WIDTH*9)         <= PriceSummaryWriter_l_inst_l_count_order_bus_wreq_addr;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid(0)                                                                <= PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid(1)                                                                <= PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid(2)                                                                <= PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid(3)                                                                <= PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid(4)                                                                <= PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid(5)                                                                <= PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid(6)                                                                <= PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid(7)                                                                <= PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid(8)                                                                <= PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_valid(9)                                                                <= PriceSummaryWriter_l_inst_l_count_order_bus_wdat_valid;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe(BUS_DATA_WIDTH/8-1 downto 0)                                     <= PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_strobe;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe(BUS_DATA_WIDTH/8+BUS_DATA_WIDTH/8-1 downto BUS_DATA_WIDTH/8)     <= PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_strobe;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe(BUS_DATA_WIDTH/8*2+BUS_DATA_WIDTH/8-1 downto BUS_DATA_WIDTH/8*2) <= PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_strobe;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe(BUS_DATA_WIDTH/8*3+BUS_DATA_WIDTH/8-1 downto BUS_DATA_WIDTH/8*3) <= PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_strobe;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe(BUS_DATA_WIDTH/8*4+BUS_DATA_WIDTH/8-1 downto BUS_DATA_WIDTH/8*4) <= PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_strobe;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe(BUS_DATA_WIDTH/8*5+BUS_DATA_WIDTH/8-1 downto BUS_DATA_WIDTH/8*5) <= PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_strobe;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe(BUS_DATA_WIDTH/8*6+BUS_DATA_WIDTH/8-1 downto BUS_DATA_WIDTH/8*6) <= PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_strobe;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe(BUS_DATA_WIDTH/8*7+BUS_DATA_WIDTH/8-1 downto BUS_DATA_WIDTH/8*7) <= PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_strobe;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe(BUS_DATA_WIDTH/8*8+BUS_DATA_WIDTH/8-1 downto BUS_DATA_WIDTH/8*8) <= PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_strobe;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_strobe(BUS_DATA_WIDTH/8*9+BUS_DATA_WIDTH/8-1 downto BUS_DATA_WIDTH/8*9) <= PriceSummaryWriter_l_inst_l_count_order_bus_wdat_strobe;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last(0)                                                                 <= PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_last;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last(1)                                                                 <= PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_last;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last(2)                                                                 <= PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_last;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last(3)                                                                 <= PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_last;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last(4)                                                                 <= PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_last;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last(5)                                                                 <= PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_last;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last(6)                                                                 <= PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_last;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last(7)                                                                 <= PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_last;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last(8)                                                                 <= PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_last;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_last(9)                                                                 <= PriceSummaryWriter_l_inst_l_count_order_bus_wdat_last;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data(BUS_DATA_WIDTH-1 downto 0)                                         <= PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_data;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data(BUS_DATA_WIDTH+BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH)             <= PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_data;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data(BUS_DATA_WIDTH*2+BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH*2)         <= PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_data;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data(BUS_DATA_WIDTH*3+BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH*3)         <= PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_data;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data(BUS_DATA_WIDTH*4+BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH*4)         <= PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_data;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data(BUS_DATA_WIDTH*5+BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH*5)         <= PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_data;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data(BUS_DATA_WIDTH*6+BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH*6)         <= PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_data;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data(BUS_DATA_WIDTH*7+BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH*7)         <= PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_data;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data(BUS_DATA_WIDTH*8+BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH*8)         <= PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_data;
  WRAW64DW512LW8BS1BM16_inst_bsv_wdat_data(BUS_DATA_WIDTH*9+BUS_DATA_WIDTH-1 downto BUS_DATA_WIDTH*9)         <= PriceSummaryWriter_l_inst_l_count_order_bus_wdat_data;
  PriceSummaryWriter_l_inst_l_sum_qty_bus_wreq_ready                                                          <= WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready(2);
  PriceSummaryWriter_l_inst_l_sum_qty_bus_wdat_ready                                                          <= WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready(2);
  PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wreq_ready                                                   <= WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready(4);
  PriceSummaryWriter_l_inst_l_sum_disc_price_bus_wdat_ready                                                   <= WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready(4);
  PriceSummaryWriter_l_inst_l_sum_charge_bus_wreq_ready                                                       <= WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready(5);
  PriceSummaryWriter_l_inst_l_sum_charge_bus_wdat_ready                                                       <= WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready(5);
  PriceSummaryWriter_l_inst_l_sum_base_price_bus_wreq_ready                                                   <= WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready(3);
  PriceSummaryWriter_l_inst_l_sum_base_price_bus_wdat_ready                                                   <= WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready(3);
  PriceSummaryWriter_l_inst_l_returnflag_o_bus_wreq_ready                                                     <= WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready(0);
  PriceSummaryWriter_l_inst_l_returnflag_o_bus_wdat_ready                                                     <= WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready(0);
  PriceSummaryWriter_l_inst_l_linestatus_o_bus_wreq_ready                                                     <= WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready(1);
  PriceSummaryWriter_l_inst_l_linestatus_o_bus_wdat_ready                                                     <= WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready(1);
  PriceSummaryWriter_l_inst_l_count_order_bus_wreq_ready                                                      <= WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready(9);
  PriceSummaryWriter_l_inst_l_count_order_bus_wdat_ready                                                      <= WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready(9);
  PriceSummaryWriter_l_inst_l_avg_qty_bus_wreq_ready                                                          <= WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready(6);
  PriceSummaryWriter_l_inst_l_avg_qty_bus_wdat_ready                                                          <= WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready(6);
  PriceSummaryWriter_l_inst_l_avg_price_bus_wreq_ready                                                        <= WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready(7);
  PriceSummaryWriter_l_inst_l_avg_price_bus_wdat_ready                                                        <= WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready(7);
  PriceSummaryWriter_l_inst_l_avg_disc_bus_wreq_ready                                                         <= WRAW64DW512LW8BS1BM16_inst_bsv_wreq_ready(8);
  PriceSummaryWriter_l_inst_l_avg_disc_bus_wdat_ready                                                         <= WRAW64DW512LW8BS1BM16_inst_bsv_wdat_ready(8);

end architecture;
