-- Copyright 2018-2019 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
-- This file was generated by Fletchgen. Modify this file at your own risk.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library work;
use work.Array_pkg.all;
use work.mmio_pkg.all;

entity PriceSummary_Nucleus is
  generic (
    INDEX_WIDTH                    : integer := 32;
    TAG_WIDTH                      : integer := 1;
    L_QUANTITY_BUS_ADDR_WIDTH      : integer := 64;
    L_EXTENDEDPRICE_BUS_ADDR_WIDTH : integer := 64;
    L_DISCOUNT_BUS_ADDR_WIDTH      : integer := 64;
    L_TAX_BUS_ADDR_WIDTH           : integer := 64;
    L_RETURNFLAG_BUS_ADDR_WIDTH    : integer := 64;
    L_LINESTATUS_BUS_ADDR_WIDTH    : integer := 64;
    L_SHIPDATE_BUS_ADDR_WIDTH      : integer := 64
  );
  port (
    kcd_clk                      : in  std_logic;
    kcd_reset                    : in  std_logic;
    mmio_awvalid                 : in  std_logic;
    mmio_awready                 : out std_logic;
    mmio_awaddr                  : in  std_logic_vector(31 downto 0);
    mmio_wvalid                  : in  std_logic;
    mmio_wready                  : out std_logic;
    mmio_wdata                   : in  std_logic_vector(31 downto 0);
    mmio_wstrb                   : in  std_logic_vector(3 downto 0);
    mmio_bvalid                  : out std_logic;
    mmio_bready                  : in  std_logic;
    mmio_bresp                   : out std_logic_vector(1 downto 0);
    mmio_arvalid                 : in  std_logic;
    mmio_arready                 : out std_logic;
    mmio_araddr                  : in  std_logic_vector(31 downto 0);
    mmio_rvalid                  : out std_logic;
    mmio_rready                  : in  std_logic;
    mmio_rdata                   : out std_logic_vector(31 downto 0);
    mmio_rresp                   : out std_logic_vector(1 downto 0);
    l_quantity_valid             : in  std_logic;
    l_quantity_ready             : out std_logic;
    l_quantity_dvalid            : in  std_logic;
    l_quantity_last              : in  std_logic;
    l_quantity                   : in  std_logic_vector(63 downto 0);
    l_extendedprice_valid        : in  std_logic;
    l_extendedprice_ready        : out std_logic;
    l_extendedprice_dvalid       : in  std_logic;
    l_extendedprice_last         : in  std_logic;
    l_extendedprice              : in  std_logic_vector(63 downto 0);
    l_discount_valid             : in  std_logic;
    l_discount_ready             : out std_logic;
    l_discount_dvalid            : in  std_logic;
    l_discount_last              : in  std_logic;
    l_discount                   : in  std_logic_vector(63 downto 0);
    l_tax_valid                  : in  std_logic;
    l_tax_ready                  : out std_logic;
    l_tax_dvalid                 : in  std_logic;
    l_tax_last                   : in  std_logic;
    l_tax                        : in  std_logic_vector(63 downto 0);
    l_returnflag_valid           : in  std_logic;
    l_returnflag_ready           : out std_logic;
    l_returnflag_dvalid          : in  std_logic;
    l_returnflag_last            : in  std_logic;
    l_returnflag_length          : in  std_logic_vector(31 downto 0);
    l_returnflag_count           : in  std_logic_vector(0 downto 0);
    l_returnflag_chars_valid     : in  std_logic;
    l_returnflag_chars_ready     : out std_logic;
    l_returnflag_chars_dvalid    : in  std_logic;
    l_returnflag_chars_last      : in  std_logic;
    l_returnflag_chars           : in  std_logic_vector(7 downto 0);
    l_returnflag_chars_count     : in  std_logic_vector(0 downto 0);
    l_linestatus_valid           : in  std_logic;
    l_linestatus_ready           : out std_logic;
    l_linestatus_dvalid          : in  std_logic;
    l_linestatus_last            : in  std_logic;
    l_linestatus_length          : in  std_logic_vector(31 downto 0);
    l_linestatus_count           : in  std_logic_vector(0 downto 0);
    l_linestatus_chars_valid     : in  std_logic;
    l_linestatus_chars_ready     : out std_logic;
    l_linestatus_chars_dvalid    : in  std_logic;
    l_linestatus_chars_last      : in  std_logic;
    l_linestatus_chars           : in  std_logic_vector(7 downto 0);
    l_linestatus_chars_count     : in  std_logic_vector(0 downto 0);
    l_shipdate_valid             : in  std_logic;
    l_shipdate_ready             : out std_logic;
    l_shipdate_dvalid            : in  std_logic;
    l_shipdate_last              : in  std_logic;
    l_shipdate                   : in  std_logic_vector(31 downto 0);
    l_quantity_unl_valid         : in  std_logic;
    l_quantity_unl_ready         : out std_logic;
    l_quantity_unl_tag           : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_extendedprice_unl_valid    : in  std_logic;
    l_extendedprice_unl_ready    : out std_logic;
    l_extendedprice_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_discount_unl_valid         : in  std_logic;
    l_discount_unl_ready         : out std_logic;
    l_discount_unl_tag           : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_tax_unl_valid              : in  std_logic;
    l_tax_unl_ready              : out std_logic;
    l_tax_unl_tag                : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_returnflag_unl_valid       : in  std_logic;
    l_returnflag_unl_ready       : out std_logic;
    l_returnflag_unl_tag         : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_linestatus_unl_valid       : in  std_logic;
    l_linestatus_unl_ready       : out std_logic;
    l_linestatus_unl_tag         : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_shipdate_unl_valid         : in  std_logic;
    l_shipdate_unl_ready         : out std_logic;
    l_shipdate_unl_tag           : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_quantity_cmd_valid         : out std_logic;
    l_quantity_cmd_ready         : in  std_logic;
    l_quantity_cmd_firstIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_quantity_cmd_lastIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_quantity_cmd_ctrl          : out std_logic_vector(L_QUANTITY_BUS_ADDR_WIDTH-1 downto 0);
    l_quantity_cmd_tag           : out std_logic_vector(TAG_WIDTH-1 downto 0);
    l_extendedprice_cmd_valid    : out std_logic;
    l_extendedprice_cmd_ready    : in  std_logic;
    l_extendedprice_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_extendedprice_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_extendedprice_cmd_ctrl     : out std_logic_vector(L_EXTENDEDPRICE_BUS_ADDR_WIDTH-1 downto 0);
    l_extendedprice_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
    l_discount_cmd_valid         : out std_logic;
    l_discount_cmd_ready         : in  std_logic;
    l_discount_cmd_firstIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_discount_cmd_lastIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_discount_cmd_ctrl          : out std_logic_vector(L_DISCOUNT_BUS_ADDR_WIDTH-1 downto 0);
    l_discount_cmd_tag           : out std_logic_vector(TAG_WIDTH-1 downto 0);
    l_tax_cmd_valid              : out std_logic;
    l_tax_cmd_ready              : in  std_logic;
    l_tax_cmd_firstIdx           : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_tax_cmd_lastIdx            : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_tax_cmd_ctrl               : out std_logic_vector(L_TAX_BUS_ADDR_WIDTH-1 downto 0);
    l_tax_cmd_tag                : out std_logic_vector(TAG_WIDTH-1 downto 0);
    l_returnflag_cmd_valid       : out std_logic;
    l_returnflag_cmd_ready       : in  std_logic;
    l_returnflag_cmd_firstIdx    : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_returnflag_cmd_lastIdx     : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_returnflag_cmd_ctrl        : out std_logic_vector(L_RETURNFLAG_BUS_ADDR_WIDTH*2-1 downto 0);
    l_returnflag_cmd_tag         : out std_logic_vector(TAG_WIDTH-1 downto 0);
    l_linestatus_cmd_valid       : out std_logic;
    l_linestatus_cmd_ready       : in  std_logic;
    l_linestatus_cmd_firstIdx    : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_linestatus_cmd_lastIdx     : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_linestatus_cmd_ctrl        : out std_logic_vector(L_LINESTATUS_BUS_ADDR_WIDTH*2-1 downto 0);
    l_linestatus_cmd_tag         : out std_logic_vector(TAG_WIDTH-1 downto 0);
    l_shipdate_cmd_valid         : out std_logic;
    l_shipdate_cmd_ready         : in  std_logic;
    l_shipdate_cmd_firstIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_shipdate_cmd_lastIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_shipdate_cmd_ctrl          : out std_logic_vector(L_SHIPDATE_BUS_ADDR_WIDTH-1 downto 0);
    l_shipdate_cmd_tag           : out std_logic_vector(TAG_WIDTH-1 downto 0)
  );
end entity;

architecture Implementation of PriceSummary_Nucleus is
  component PriceSummary is
    generic (
      INDEX_WIDTH : integer := 32;
      TAG_WIDTH   : integer := 1
    );
    port (
      kcd_clk                      : in  std_logic;
      kcd_reset                    : in  std_logic;
      l_quantity_valid             : in  std_logic;
      l_quantity_ready             : out std_logic;
      l_quantity_dvalid            : in  std_logic;
      l_quantity_last              : in  std_logic;
      l_quantity                   : in  std_logic_vector(63 downto 0);
      l_extendedprice_valid        : in  std_logic;
      l_extendedprice_ready        : out std_logic;
      l_extendedprice_dvalid       : in  std_logic;
      l_extendedprice_last         : in  std_logic;
      l_extendedprice              : in  std_logic_vector(63 downto 0);
      l_discount_valid             : in  std_logic;
      l_discount_ready             : out std_logic;
      l_discount_dvalid            : in  std_logic;
      l_discount_last              : in  std_logic;
      l_discount                   : in  std_logic_vector(63 downto 0);
      l_tax_valid                  : in  std_logic;
      l_tax_ready                  : out std_logic;
      l_tax_dvalid                 : in  std_logic;
      l_tax_last                   : in  std_logic;
      l_tax                        : in  std_logic_vector(63 downto 0);
      l_returnflag_valid           : in  std_logic;
      l_returnflag_ready           : out std_logic;
      l_returnflag_dvalid          : in  std_logic;
      l_returnflag_last            : in  std_logic;
      l_returnflag_length          : in  std_logic_vector(31 downto 0);
      l_returnflag_count           : in  std_logic_vector(0 downto 0);
      l_returnflag_chars_valid     : in  std_logic;
      l_returnflag_chars_ready     : out std_logic;
      l_returnflag_chars_dvalid    : in  std_logic;
      l_returnflag_chars_last      : in  std_logic;
      l_returnflag_chars           : in  std_logic_vector(7 downto 0);
      l_returnflag_chars_count     : in  std_logic_vector(0 downto 0);
      l_linestatus_valid           : in  std_logic;
      l_linestatus_ready           : out std_logic;
      l_linestatus_dvalid          : in  std_logic;
      l_linestatus_last            : in  std_logic;
      l_linestatus_length          : in  std_logic_vector(31 downto 0);
      l_linestatus_count           : in  std_logic_vector(0 downto 0);
      l_linestatus_chars_valid     : in  std_logic;
      l_linestatus_chars_ready     : out std_logic;
      l_linestatus_chars_dvalid    : in  std_logic;
      l_linestatus_chars_last      : in  std_logic;
      l_linestatus_chars           : in  std_logic_vector(7 downto 0);
      l_linestatus_chars_count     : in  std_logic_vector(0 downto 0);
      l_shipdate_valid             : in  std_logic;
      l_shipdate_ready             : out std_logic;
      l_shipdate_dvalid            : in  std_logic;
      l_shipdate_last              : in  std_logic;
      l_shipdate                   : in  std_logic_vector(31 downto 0);
      l_quantity_unl_valid         : in  std_logic;
      l_quantity_unl_ready         : out std_logic;
      l_quantity_unl_tag           : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_extendedprice_unl_valid    : in  std_logic;
      l_extendedprice_unl_ready    : out std_logic;
      l_extendedprice_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_discount_unl_valid         : in  std_logic;
      l_discount_unl_ready         : out std_logic;
      l_discount_unl_tag           : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_tax_unl_valid              : in  std_logic;
      l_tax_unl_ready              : out std_logic;
      l_tax_unl_tag                : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_returnflag_unl_valid       : in  std_logic;
      l_returnflag_unl_ready       : out std_logic;
      l_returnflag_unl_tag         : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_linestatus_unl_valid       : in  std_logic;
      l_linestatus_unl_ready       : out std_logic;
      l_linestatus_unl_tag         : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_shipdate_unl_valid         : in  std_logic;
      l_shipdate_unl_ready         : out std_logic;
      l_shipdate_unl_tag           : in  std_logic_vector(TAG_WIDTH-1 downto 0);
      l_quantity_cmd_valid         : out std_logic;
      l_quantity_cmd_ready         : in  std_logic;
      l_quantity_cmd_firstIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_quantity_cmd_lastIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_quantity_cmd_tag           : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_extendedprice_cmd_valid    : out std_logic;
      l_extendedprice_cmd_ready    : in  std_logic;
      l_extendedprice_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_extendedprice_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_extendedprice_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_discount_cmd_valid         : out std_logic;
      l_discount_cmd_ready         : in  std_logic;
      l_discount_cmd_firstIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_discount_cmd_lastIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_discount_cmd_tag           : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_tax_cmd_valid              : out std_logic;
      l_tax_cmd_ready              : in  std_logic;
      l_tax_cmd_firstIdx           : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_tax_cmd_lastIdx            : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_tax_cmd_tag                : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_returnflag_cmd_valid       : out std_logic;
      l_returnflag_cmd_ready       : in  std_logic;
      l_returnflag_cmd_firstIdx    : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_returnflag_cmd_lastIdx     : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_returnflag_cmd_tag         : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_linestatus_cmd_valid       : out std_logic;
      l_linestatus_cmd_ready       : in  std_logic;
      l_linestatus_cmd_firstIdx    : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_linestatus_cmd_lastIdx     : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_linestatus_cmd_tag         : out std_logic_vector(TAG_WIDTH-1 downto 0);
      l_shipdate_cmd_valid         : out std_logic;
      l_shipdate_cmd_ready         : in  std_logic;
      l_shipdate_cmd_firstIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_shipdate_cmd_lastIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
      l_shipdate_cmd_tag           : out std_logic_vector(TAG_WIDTH-1 downto 0);
      start                        : in  std_logic;
      stop                         : in  std_logic;
      reset                        : in  std_logic;
      idle                         : out std_logic;
      busy                         : out std_logic;
      done                         : out std_logic;
      result                       : out std_logic_vector(63 downto 0);
      l_firstidx                   : in  std_logic_vector(31 downto 0);
      l_lastidx                    : in  std_logic_vector(31 downto 0);
      rhigh                        : out std_logic_vector(31 downto 0);
      rlow                         : out std_logic_vector(31 downto 0);
      status_1                     : out std_logic_vector(31 downto 0);
      status_2                     : out std_logic_vector(31 downto 0);
      r1                           : out std_logic_vector(63 downto 0);
      r2                           : out std_logic_vector(63 downto 0);
      r3                           : out std_logic_vector(63 downto 0);
      r4                           : out std_logic_vector(63 downto 0);
      r5                           : out std_logic_vector(63 downto 0);
      r6                           : out std_logic_vector(63 downto 0);
      r7                           : out std_logic_vector(63 downto 0);
      r8                           : out std_logic_vector(63 downto 0)
    );
  end component;

  signal PriceSummary_inst_l_quantity_valid                 : std_logic;
  signal PriceSummary_inst_l_quantity_ready                 : std_logic;
  signal PriceSummary_inst_l_quantity_dvalid                : std_logic;
  signal PriceSummary_inst_l_quantity_last                  : std_logic;
  signal PriceSummary_inst_l_quantity                       : std_logic_vector(63 downto 0);

  signal PriceSummary_inst_l_extendedprice_valid            : std_logic;
  signal PriceSummary_inst_l_extendedprice_ready            : std_logic;
  signal PriceSummary_inst_l_extendedprice_dvalid           : std_logic;
  signal PriceSummary_inst_l_extendedprice_last             : std_logic;
  signal PriceSummary_inst_l_extendedprice                  : std_logic_vector(63 downto 0);

  signal PriceSummary_inst_l_discount_valid                 : std_logic;
  signal PriceSummary_inst_l_discount_ready                 : std_logic;
  signal PriceSummary_inst_l_discount_dvalid                : std_logic;
  signal PriceSummary_inst_l_discount_last                  : std_logic;
  signal PriceSummary_inst_l_discount                       : std_logic_vector(63 downto 0);

  signal PriceSummary_inst_l_tax_valid                      : std_logic;
  signal PriceSummary_inst_l_tax_ready                      : std_logic;
  signal PriceSummary_inst_l_tax_dvalid                     : std_logic;
  signal PriceSummary_inst_l_tax_last                       : std_logic;
  signal PriceSummary_inst_l_tax                            : std_logic_vector(63 downto 0);

  signal PriceSummary_inst_l_returnflag_valid               : std_logic;
  signal PriceSummary_inst_l_returnflag_ready               : std_logic;
  signal PriceSummary_inst_l_returnflag_dvalid              : std_logic;
  signal PriceSummary_inst_l_returnflag_last                : std_logic;
  signal PriceSummary_inst_l_returnflag_length              : std_logic_vector(31 downto 0);
  signal PriceSummary_inst_l_returnflag_count               : std_logic_vector(0 downto 0);
  signal PriceSummary_inst_l_returnflag_chars_valid         : std_logic;
  signal PriceSummary_inst_l_returnflag_chars_ready         : std_logic;
  signal PriceSummary_inst_l_returnflag_chars_dvalid        : std_logic;
  signal PriceSummary_inst_l_returnflag_chars_last          : std_logic;
  signal PriceSummary_inst_l_returnflag_chars               : std_logic_vector(7 downto 0);
  signal PriceSummary_inst_l_returnflag_chars_count         : std_logic_vector(0 downto 0);

  signal PriceSummary_inst_l_linestatus_valid               : std_logic;
  signal PriceSummary_inst_l_linestatus_ready               : std_logic;
  signal PriceSummary_inst_l_linestatus_dvalid              : std_logic;
  signal PriceSummary_inst_l_linestatus_last                : std_logic;
  signal PriceSummary_inst_l_linestatus_length              : std_logic_vector(31 downto 0);
  signal PriceSummary_inst_l_linestatus_count               : std_logic_vector(0 downto 0);
  signal PriceSummary_inst_l_linestatus_chars_valid         : std_logic;
  signal PriceSummary_inst_l_linestatus_chars_ready         : std_logic;
  signal PriceSummary_inst_l_linestatus_chars_dvalid        : std_logic;
  signal PriceSummary_inst_l_linestatus_chars_last          : std_logic;
  signal PriceSummary_inst_l_linestatus_chars               : std_logic_vector(7 downto 0);
  signal PriceSummary_inst_l_linestatus_chars_count         : std_logic_vector(0 downto 0);

  signal PriceSummary_inst_l_shipdate_valid                 : std_logic;
  signal PriceSummary_inst_l_shipdate_ready                 : std_logic;
  signal PriceSummary_inst_l_shipdate_dvalid                : std_logic;
  signal PriceSummary_inst_l_shipdate_last                  : std_logic;
  signal PriceSummary_inst_l_shipdate                       : std_logic_vector(31 downto 0);

  signal PriceSummary_inst_l_quantity_unl_valid             : std_logic;
  signal PriceSummary_inst_l_quantity_unl_ready             : std_logic;
  signal PriceSummary_inst_l_quantity_unl_tag               : std_logic_vector(0 downto 0);

  signal PriceSummary_inst_l_extendedprice_unl_valid        : std_logic;
  signal PriceSummary_inst_l_extendedprice_unl_ready        : std_logic;
  signal PriceSummary_inst_l_extendedprice_unl_tag          : std_logic_vector(0 downto 0);

  signal PriceSummary_inst_l_discount_unl_valid             : std_logic;
  signal PriceSummary_inst_l_discount_unl_ready             : std_logic;
  signal PriceSummary_inst_l_discount_unl_tag               : std_logic_vector(0 downto 0);

  signal PriceSummary_inst_l_tax_unl_valid                  : std_logic;
  signal PriceSummary_inst_l_tax_unl_ready                  : std_logic;
  signal PriceSummary_inst_l_tax_unl_tag                    : std_logic_vector(0 downto 0);

  signal PriceSummary_inst_l_returnflag_unl_valid           : std_logic;
  signal PriceSummary_inst_l_returnflag_unl_ready           : std_logic;
  signal PriceSummary_inst_l_returnflag_unl_tag             : std_logic_vector(0 downto 0);

  signal PriceSummary_inst_l_linestatus_unl_valid           : std_logic;
  signal PriceSummary_inst_l_linestatus_unl_ready           : std_logic;
  signal PriceSummary_inst_l_linestatus_unl_tag             : std_logic_vector(0 downto 0);

  signal PriceSummary_inst_l_shipdate_unl_valid             : std_logic;
  signal PriceSummary_inst_l_shipdate_unl_ready             : std_logic;
  signal PriceSummary_inst_l_shipdate_unl_tag               : std_logic_vector(0 downto 0);

  signal PriceSummary_inst_l_quantity_cmd_valid             : std_logic;
  signal PriceSummary_inst_l_quantity_cmd_ready             : std_logic;
  signal PriceSummary_inst_l_quantity_cmd_firstIdx          : std_logic_vector(31 downto 0);
  signal PriceSummary_inst_l_quantity_cmd_lastIdx           : std_logic_vector(31 downto 0);
  signal PriceSummary_inst_l_quantity_cmd_tag               : std_logic_vector(0 downto 0);

  signal PriceSummary_inst_l_extendedprice_cmd_valid        : std_logic;
  signal PriceSummary_inst_l_extendedprice_cmd_ready        : std_logic;
  signal PriceSummary_inst_l_extendedprice_cmd_firstIdx     : std_logic_vector(31 downto 0);
  signal PriceSummary_inst_l_extendedprice_cmd_lastIdx      : std_logic_vector(31 downto 0);
  signal PriceSummary_inst_l_extendedprice_cmd_tag          : std_logic_vector(0 downto 0);

  signal PriceSummary_inst_l_discount_cmd_valid             : std_logic;
  signal PriceSummary_inst_l_discount_cmd_ready             : std_logic;
  signal PriceSummary_inst_l_discount_cmd_firstIdx          : std_logic_vector(31 downto 0);
  signal PriceSummary_inst_l_discount_cmd_lastIdx           : std_logic_vector(31 downto 0);
  signal PriceSummary_inst_l_discount_cmd_tag               : std_logic_vector(0 downto 0);

  signal PriceSummary_inst_l_tax_cmd_valid                  : std_logic;
  signal PriceSummary_inst_l_tax_cmd_ready                  : std_logic;
  signal PriceSummary_inst_l_tax_cmd_firstIdx               : std_logic_vector(31 downto 0);
  signal PriceSummary_inst_l_tax_cmd_lastIdx                : std_logic_vector(31 downto 0);
  signal PriceSummary_inst_l_tax_cmd_tag                    : std_logic_vector(0 downto 0);

  signal PriceSummary_inst_l_returnflag_cmd_valid           : std_logic;
  signal PriceSummary_inst_l_returnflag_cmd_ready           : std_logic;
  signal PriceSummary_inst_l_returnflag_cmd_firstIdx        : std_logic_vector(31 downto 0);
  signal PriceSummary_inst_l_returnflag_cmd_lastIdx         : std_logic_vector(31 downto 0);
  signal PriceSummary_inst_l_returnflag_cmd_tag             : std_logic_vector(0 downto 0);

  signal PriceSummary_inst_l_linestatus_cmd_valid           : std_logic;
  signal PriceSummary_inst_l_linestatus_cmd_ready           : std_logic;
  signal PriceSummary_inst_l_linestatus_cmd_firstIdx        : std_logic_vector(31 downto 0);
  signal PriceSummary_inst_l_linestatus_cmd_lastIdx         : std_logic_vector(31 downto 0);
  signal PriceSummary_inst_l_linestatus_cmd_tag             : std_logic_vector(0 downto 0);

  signal PriceSummary_inst_l_shipdate_cmd_valid             : std_logic;
  signal PriceSummary_inst_l_shipdate_cmd_ready             : std_logic;
  signal PriceSummary_inst_l_shipdate_cmd_firstIdx          : std_logic_vector(31 downto 0);
  signal PriceSummary_inst_l_shipdate_cmd_lastIdx           : std_logic_vector(31 downto 0);
  signal PriceSummary_inst_l_shipdate_cmd_tag               : std_logic_vector(0 downto 0);

  signal PriceSummary_inst_start                            : std_logic;
  signal PriceSummary_inst_stop                             : std_logic;
  signal PriceSummary_inst_reset                            : std_logic;
  signal PriceSummary_inst_idle                             : std_logic;
  signal PriceSummary_inst_busy                             : std_logic;
  signal PriceSummary_inst_done                             : std_logic;
  signal PriceSummary_inst_result                           : std_logic_vector(63 downto 0);
  signal PriceSummary_inst_l_firstidx                       : std_logic_vector(31 downto 0);
  signal PriceSummary_inst_l_lastidx                        : std_logic_vector(31 downto 0);
  signal PriceSummary_inst_rhigh                            : std_logic_vector(31 downto 0);
  signal PriceSummary_inst_rlow                             : std_logic_vector(31 downto 0);
  signal PriceSummary_inst_status_1                         : std_logic_vector(31 downto 0);
  signal PriceSummary_inst_status_2                         : std_logic_vector(31 downto 0);
  signal PriceSummary_inst_r1                               : std_logic_vector(63 downto 0);
  signal PriceSummary_inst_r2                               : std_logic_vector(63 downto 0);
  signal PriceSummary_inst_r3                               : std_logic_vector(63 downto 0);
  signal PriceSummary_inst_r4                               : std_logic_vector(63 downto 0);
  signal PriceSummary_inst_r5                               : std_logic_vector(63 downto 0);
  signal PriceSummary_inst_r6                               : std_logic_vector(63 downto 0);
  signal PriceSummary_inst_r7                               : std_logic_vector(63 downto 0);
  signal PriceSummary_inst_r8                               : std_logic_vector(63 downto 0);
  signal mmio_inst_f_start_data                             : std_logic;
  signal mmio_inst_f_stop_data                              : std_logic;
  signal mmio_inst_f_reset_data                             : std_logic;
  signal mmio_inst_f_idle_write_data                        : std_logic;
  signal mmio_inst_f_busy_write_data                        : std_logic;
  signal mmio_inst_f_done_write_data                        : std_logic;
  signal mmio_inst_f_result_write_data                      : std_logic_vector(63 downto 0);
  signal mmio_inst_f_l_firstidx_data                        : std_logic_vector(31 downto 0);
  signal mmio_inst_f_l_lastidx_data                         : std_logic_vector(31 downto 0);
  signal mmio_inst_f_l_quantity_values_data                 : std_logic_vector(63 downto 0);
  signal mmio_inst_f_l_extendedprice_values_data            : std_logic_vector(63 downto 0);
  signal mmio_inst_f_l_discount_values_data                 : std_logic_vector(63 downto 0);
  signal mmio_inst_f_l_tax_values_data                      : std_logic_vector(63 downto 0);
  signal mmio_inst_f_l_returnflag_offsets_data              : std_logic_vector(63 downto 0);
  signal mmio_inst_f_l_returnflag_values_data               : std_logic_vector(63 downto 0);
  signal mmio_inst_f_l_linestatus_offsets_data              : std_logic_vector(63 downto 0);
  signal mmio_inst_f_l_linestatus_values_data               : std_logic_vector(63 downto 0);
  signal mmio_inst_f_l_shipdate_values_data                 : std_logic_vector(63 downto 0);
  signal mmio_inst_f_rhigh_write_data                       : std_logic_vector(31 downto 0);
  signal mmio_inst_f_rlow_write_data                        : std_logic_vector(31 downto 0);
  signal mmio_inst_f_status_1_write_data                    : std_logic_vector(31 downto 0);
  signal mmio_inst_f_status_2_write_data                    : std_logic_vector(31 downto 0);
  signal mmio_inst_f_r1_write_data                          : std_logic_vector(63 downto 0);
  signal mmio_inst_f_r2_write_data                          : std_logic_vector(63 downto 0);
  signal mmio_inst_f_r3_write_data                          : std_logic_vector(63 downto 0);
  signal mmio_inst_f_r4_write_data                          : std_logic_vector(63 downto 0);
  signal mmio_inst_f_r5_write_data                          : std_logic_vector(63 downto 0);
  signal mmio_inst_f_r6_write_data                          : std_logic_vector(63 downto 0);
  signal mmio_inst_f_r7_write_data                          : std_logic_vector(63 downto 0);
  signal mmio_inst_f_r8_write_data                          : std_logic_vector(63 downto 0);
  signal mmio_inst_f_Profile_enable_data                    : std_logic;
  signal mmio_inst_f_Profile_clear_data                     : std_logic;
  signal mmio_inst_mmio_awvalid                             : std_logic;
  signal mmio_inst_mmio_awready                             : std_logic;
  signal mmio_inst_mmio_awaddr                              : std_logic_vector(31 downto 0);
  signal mmio_inst_mmio_wvalid                              : std_logic;
  signal mmio_inst_mmio_wready                              : std_logic;
  signal mmio_inst_mmio_wdata                               : std_logic_vector(31 downto 0);
  signal mmio_inst_mmio_wstrb                               : std_logic_vector(3 downto 0);
  signal mmio_inst_mmio_bvalid                              : std_logic;
  signal mmio_inst_mmio_bready                              : std_logic;
  signal mmio_inst_mmio_bresp                               : std_logic_vector(1 downto 0);
  signal mmio_inst_mmio_arvalid                             : std_logic;
  signal mmio_inst_mmio_arready                             : std_logic;
  signal mmio_inst_mmio_araddr                              : std_logic_vector(31 downto 0);
  signal mmio_inst_mmio_rvalid                              : std_logic;
  signal mmio_inst_mmio_rready                              : std_logic;
  signal mmio_inst_mmio_rdata                               : std_logic_vector(31 downto 0);
  signal mmio_inst_mmio_rresp                               : std_logic_vector(1 downto 0);

  signal l_quantity_cmd_accm_inst_kernel_cmd_valid          : std_logic;
  signal l_quantity_cmd_accm_inst_kernel_cmd_ready          : std_logic;
  signal l_quantity_cmd_accm_inst_kernel_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_quantity_cmd_accm_inst_kernel_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_quantity_cmd_accm_inst_kernel_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_quantity_cmd_accm_inst_nucleus_cmd_valid         : std_logic;
  signal l_quantity_cmd_accm_inst_nucleus_cmd_ready         : std_logic;
  signal l_quantity_cmd_accm_inst_nucleus_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_quantity_cmd_accm_inst_nucleus_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_quantity_cmd_accm_inst_nucleus_cmd_ctrl          : std_logic_vector(L_QUANTITY_BUS_ADDR_WIDTH-1 downto 0);
  signal l_quantity_cmd_accm_inst_nucleus_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_extendedprice_cmd_accm_inst_kernel_cmd_valid     : std_logic;
  signal l_extendedprice_cmd_accm_inst_kernel_cmd_ready     : std_logic;
  signal l_extendedprice_cmd_accm_inst_kernel_cmd_firstIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_extendedprice_cmd_accm_inst_kernel_cmd_lastIdx   : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_extendedprice_cmd_accm_inst_kernel_cmd_tag       : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_extendedprice_cmd_accm_inst_nucleus_cmd_valid    : std_logic;
  signal l_extendedprice_cmd_accm_inst_nucleus_cmd_ready    : std_logic;
  signal l_extendedprice_cmd_accm_inst_nucleus_cmd_firstIdx : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_extendedprice_cmd_accm_inst_nucleus_cmd_lastIdx  : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_extendedprice_cmd_accm_inst_nucleus_cmd_ctrl     : std_logic_vector(L_EXTENDEDPRICE_BUS_ADDR_WIDTH-1 downto 0);
  signal l_extendedprice_cmd_accm_inst_nucleus_cmd_tag      : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_discount_cmd_accm_inst_kernel_cmd_valid          : std_logic;
  signal l_discount_cmd_accm_inst_kernel_cmd_ready          : std_logic;
  signal l_discount_cmd_accm_inst_kernel_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_discount_cmd_accm_inst_kernel_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_discount_cmd_accm_inst_kernel_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_discount_cmd_accm_inst_nucleus_cmd_valid         : std_logic;
  signal l_discount_cmd_accm_inst_nucleus_cmd_ready         : std_logic;
  signal l_discount_cmd_accm_inst_nucleus_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_discount_cmd_accm_inst_nucleus_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_discount_cmd_accm_inst_nucleus_cmd_ctrl          : std_logic_vector(L_DISCOUNT_BUS_ADDR_WIDTH-1 downto 0);
  signal l_discount_cmd_accm_inst_nucleus_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_tax_cmd_accm_inst_kernel_cmd_valid               : std_logic;
  signal l_tax_cmd_accm_inst_kernel_cmd_ready               : std_logic;
  signal l_tax_cmd_accm_inst_kernel_cmd_firstIdx            : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_tax_cmd_accm_inst_kernel_cmd_lastIdx             : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_tax_cmd_accm_inst_kernel_cmd_tag                 : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_tax_cmd_accm_inst_nucleus_cmd_valid              : std_logic;
  signal l_tax_cmd_accm_inst_nucleus_cmd_ready              : std_logic;
  signal l_tax_cmd_accm_inst_nucleus_cmd_firstIdx           : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_tax_cmd_accm_inst_nucleus_cmd_lastIdx            : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_tax_cmd_accm_inst_nucleus_cmd_ctrl               : std_logic_vector(L_TAX_BUS_ADDR_WIDTH-1 downto 0);
  signal l_tax_cmd_accm_inst_nucleus_cmd_tag                : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_returnflag_cmd_accm_inst_kernel_cmd_valid        : std_logic;
  signal l_returnflag_cmd_accm_inst_kernel_cmd_ready        : std_logic;
  signal l_returnflag_cmd_accm_inst_kernel_cmd_firstIdx     : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_returnflag_cmd_accm_inst_kernel_cmd_lastIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_returnflag_cmd_accm_inst_kernel_cmd_tag          : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_returnflag_cmd_accm_inst_nucleus_cmd_valid       : std_logic;
  signal l_returnflag_cmd_accm_inst_nucleus_cmd_ready       : std_logic;
  signal l_returnflag_cmd_accm_inst_nucleus_cmd_firstIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_returnflag_cmd_accm_inst_nucleus_cmd_lastIdx     : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_returnflag_cmd_accm_inst_nucleus_cmd_ctrl        : std_logic_vector(2*L_RETURNFLAG_BUS_ADDR_WIDTH-1 downto 0);
  signal l_returnflag_cmd_accm_inst_nucleus_cmd_tag         : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_linestatus_cmd_accm_inst_kernel_cmd_valid        : std_logic;
  signal l_linestatus_cmd_accm_inst_kernel_cmd_ready        : std_logic;
  signal l_linestatus_cmd_accm_inst_kernel_cmd_firstIdx     : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_linestatus_cmd_accm_inst_kernel_cmd_lastIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_linestatus_cmd_accm_inst_kernel_cmd_tag          : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_linestatus_cmd_accm_inst_nucleus_cmd_valid       : std_logic;
  signal l_linestatus_cmd_accm_inst_nucleus_cmd_ready       : std_logic;
  signal l_linestatus_cmd_accm_inst_nucleus_cmd_firstIdx    : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_linestatus_cmd_accm_inst_nucleus_cmd_lastIdx     : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_linestatus_cmd_accm_inst_nucleus_cmd_ctrl        : std_logic_vector(2*L_LINESTATUS_BUS_ADDR_WIDTH-1 downto 0);
  signal l_linestatus_cmd_accm_inst_nucleus_cmd_tag         : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_shipdate_cmd_accm_inst_kernel_cmd_valid          : std_logic;
  signal l_shipdate_cmd_accm_inst_kernel_cmd_ready          : std_logic;
  signal l_shipdate_cmd_accm_inst_kernel_cmd_firstIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_shipdate_cmd_accm_inst_kernel_cmd_lastIdx        : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_shipdate_cmd_accm_inst_kernel_cmd_tag            : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_shipdate_cmd_accm_inst_nucleus_cmd_valid         : std_logic;
  signal l_shipdate_cmd_accm_inst_nucleus_cmd_ready         : std_logic;
  signal l_shipdate_cmd_accm_inst_nucleus_cmd_firstIdx      : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_shipdate_cmd_accm_inst_nucleus_cmd_lastIdx       : std_logic_vector(INDEX_WIDTH-1 downto 0);
  signal l_shipdate_cmd_accm_inst_nucleus_cmd_ctrl          : std_logic_vector(L_SHIPDATE_BUS_ADDR_WIDTH-1 downto 0);
  signal l_shipdate_cmd_accm_inst_nucleus_cmd_tag           : std_logic_vector(TAG_WIDTH-1 downto 0);

  signal l_quantity_cmd_accm_inst_ctrl      : std_logic_vector(L_QUANTITY_BUS_ADDR_WIDTH-1 downto 0);
  signal l_extendedprice_cmd_accm_inst_ctrl : std_logic_vector(L_EXTENDEDPRICE_BUS_ADDR_WIDTH-1 downto 0);
  signal l_discount_cmd_accm_inst_ctrl      : std_logic_vector(L_DISCOUNT_BUS_ADDR_WIDTH-1 downto 0);
  signal l_tax_cmd_accm_inst_ctrl           : std_logic_vector(L_TAX_BUS_ADDR_WIDTH-1 downto 0);
  signal l_returnflag_cmd_accm_inst_ctrl    : std_logic_vector(2*L_RETURNFLAG_BUS_ADDR_WIDTH-1 downto 0);
  signal l_linestatus_cmd_accm_inst_ctrl    : std_logic_vector(2*L_LINESTATUS_BUS_ADDR_WIDTH-1 downto 0);
  signal l_shipdate_cmd_accm_inst_ctrl      : std_logic_vector(L_SHIPDATE_BUS_ADDR_WIDTH-1 downto 0);

begin
  PriceSummary_inst : PriceSummary
    generic map (
      INDEX_WIDTH => 32,
      TAG_WIDTH   => 1
    )
    port map (
      kcd_clk                      => kcd_clk,
      kcd_reset                    => kcd_reset,
      l_quantity_valid             => PriceSummary_inst_l_quantity_valid,
      l_quantity_ready             => PriceSummary_inst_l_quantity_ready,
      l_quantity_dvalid            => PriceSummary_inst_l_quantity_dvalid,
      l_quantity_last              => PriceSummary_inst_l_quantity_last,
      l_quantity                   => PriceSummary_inst_l_quantity,
      l_extendedprice_valid        => PriceSummary_inst_l_extendedprice_valid,
      l_extendedprice_ready        => PriceSummary_inst_l_extendedprice_ready,
      l_extendedprice_dvalid       => PriceSummary_inst_l_extendedprice_dvalid,
      l_extendedprice_last         => PriceSummary_inst_l_extendedprice_last,
      l_extendedprice              => PriceSummary_inst_l_extendedprice,
      l_discount_valid             => PriceSummary_inst_l_discount_valid,
      l_discount_ready             => PriceSummary_inst_l_discount_ready,
      l_discount_dvalid            => PriceSummary_inst_l_discount_dvalid,
      l_discount_last              => PriceSummary_inst_l_discount_last,
      l_discount                   => PriceSummary_inst_l_discount,
      l_tax_valid                  => PriceSummary_inst_l_tax_valid,
      l_tax_ready                  => PriceSummary_inst_l_tax_ready,
      l_tax_dvalid                 => PriceSummary_inst_l_tax_dvalid,
      l_tax_last                   => PriceSummary_inst_l_tax_last,
      l_tax                        => PriceSummary_inst_l_tax,
      l_returnflag_valid           => PriceSummary_inst_l_returnflag_valid,
      l_returnflag_ready           => PriceSummary_inst_l_returnflag_ready,
      l_returnflag_dvalid          => PriceSummary_inst_l_returnflag_dvalid,
      l_returnflag_last            => PriceSummary_inst_l_returnflag_last,
      l_returnflag_length          => PriceSummary_inst_l_returnflag_length,
      l_returnflag_count           => PriceSummary_inst_l_returnflag_count,
      l_returnflag_chars_valid     => PriceSummary_inst_l_returnflag_chars_valid,
      l_returnflag_chars_ready     => PriceSummary_inst_l_returnflag_chars_ready,
      l_returnflag_chars_dvalid    => PriceSummary_inst_l_returnflag_chars_dvalid,
      l_returnflag_chars_last      => PriceSummary_inst_l_returnflag_chars_last,
      l_returnflag_chars           => PriceSummary_inst_l_returnflag_chars,
      l_returnflag_chars_count     => PriceSummary_inst_l_returnflag_chars_count,
      l_linestatus_valid           => PriceSummary_inst_l_linestatus_valid,
      l_linestatus_ready           => PriceSummary_inst_l_linestatus_ready,
      l_linestatus_dvalid          => PriceSummary_inst_l_linestatus_dvalid,
      l_linestatus_last            => PriceSummary_inst_l_linestatus_last,
      l_linestatus_length          => PriceSummary_inst_l_linestatus_length,
      l_linestatus_count           => PriceSummary_inst_l_linestatus_count,
      l_linestatus_chars_valid     => PriceSummary_inst_l_linestatus_chars_valid,
      l_linestatus_chars_ready     => PriceSummary_inst_l_linestatus_chars_ready,
      l_linestatus_chars_dvalid    => PriceSummary_inst_l_linestatus_chars_dvalid,
      l_linestatus_chars_last      => PriceSummary_inst_l_linestatus_chars_last,
      l_linestatus_chars           => PriceSummary_inst_l_linestatus_chars,
      l_linestatus_chars_count     => PriceSummary_inst_l_linestatus_chars_count,
      l_shipdate_valid             => PriceSummary_inst_l_shipdate_valid,
      l_shipdate_ready             => PriceSummary_inst_l_shipdate_ready,
      l_shipdate_dvalid            => PriceSummary_inst_l_shipdate_dvalid,
      l_shipdate_last              => PriceSummary_inst_l_shipdate_last,
      l_shipdate                   => PriceSummary_inst_l_shipdate,
      l_quantity_unl_valid         => PriceSummary_inst_l_quantity_unl_valid,
      l_quantity_unl_ready         => PriceSummary_inst_l_quantity_unl_ready,
      l_quantity_unl_tag           => PriceSummary_inst_l_quantity_unl_tag,
      l_extendedprice_unl_valid    => PriceSummary_inst_l_extendedprice_unl_valid,
      l_extendedprice_unl_ready    => PriceSummary_inst_l_extendedprice_unl_ready,
      l_extendedprice_unl_tag      => PriceSummary_inst_l_extendedprice_unl_tag,
      l_discount_unl_valid         => PriceSummary_inst_l_discount_unl_valid,
      l_discount_unl_ready         => PriceSummary_inst_l_discount_unl_ready,
      l_discount_unl_tag           => PriceSummary_inst_l_discount_unl_tag,
      l_tax_unl_valid              => PriceSummary_inst_l_tax_unl_valid,
      l_tax_unl_ready              => PriceSummary_inst_l_tax_unl_ready,
      l_tax_unl_tag                => PriceSummary_inst_l_tax_unl_tag,
      l_returnflag_unl_valid       => PriceSummary_inst_l_returnflag_unl_valid,
      l_returnflag_unl_ready       => PriceSummary_inst_l_returnflag_unl_ready,
      l_returnflag_unl_tag         => PriceSummary_inst_l_returnflag_unl_tag,
      l_linestatus_unl_valid       => PriceSummary_inst_l_linestatus_unl_valid,
      l_linestatus_unl_ready       => PriceSummary_inst_l_linestatus_unl_ready,
      l_linestatus_unl_tag         => PriceSummary_inst_l_linestatus_unl_tag,
      l_shipdate_unl_valid         => PriceSummary_inst_l_shipdate_unl_valid,
      l_shipdate_unl_ready         => PriceSummary_inst_l_shipdate_unl_ready,
      l_shipdate_unl_tag           => PriceSummary_inst_l_shipdate_unl_tag,
      l_quantity_cmd_valid         => PriceSummary_inst_l_quantity_cmd_valid,
      l_quantity_cmd_ready         => PriceSummary_inst_l_quantity_cmd_ready,
      l_quantity_cmd_firstIdx      => PriceSummary_inst_l_quantity_cmd_firstIdx,
      l_quantity_cmd_lastIdx       => PriceSummary_inst_l_quantity_cmd_lastIdx,
      l_quantity_cmd_tag           => PriceSummary_inst_l_quantity_cmd_tag,
      l_extendedprice_cmd_valid    => PriceSummary_inst_l_extendedprice_cmd_valid,
      l_extendedprice_cmd_ready    => PriceSummary_inst_l_extendedprice_cmd_ready,
      l_extendedprice_cmd_firstIdx => PriceSummary_inst_l_extendedprice_cmd_firstIdx,
      l_extendedprice_cmd_lastIdx  => PriceSummary_inst_l_extendedprice_cmd_lastIdx,
      l_extendedprice_cmd_tag      => PriceSummary_inst_l_extendedprice_cmd_tag,
      l_discount_cmd_valid         => PriceSummary_inst_l_discount_cmd_valid,
      l_discount_cmd_ready         => PriceSummary_inst_l_discount_cmd_ready,
      l_discount_cmd_firstIdx      => PriceSummary_inst_l_discount_cmd_firstIdx,
      l_discount_cmd_lastIdx       => PriceSummary_inst_l_discount_cmd_lastIdx,
      l_discount_cmd_tag           => PriceSummary_inst_l_discount_cmd_tag,
      l_tax_cmd_valid              => PriceSummary_inst_l_tax_cmd_valid,
      l_tax_cmd_ready              => PriceSummary_inst_l_tax_cmd_ready,
      l_tax_cmd_firstIdx           => PriceSummary_inst_l_tax_cmd_firstIdx,
      l_tax_cmd_lastIdx            => PriceSummary_inst_l_tax_cmd_lastIdx,
      l_tax_cmd_tag                => PriceSummary_inst_l_tax_cmd_tag,
      l_returnflag_cmd_valid       => PriceSummary_inst_l_returnflag_cmd_valid,
      l_returnflag_cmd_ready       => PriceSummary_inst_l_returnflag_cmd_ready,
      l_returnflag_cmd_firstIdx    => PriceSummary_inst_l_returnflag_cmd_firstIdx,
      l_returnflag_cmd_lastIdx     => PriceSummary_inst_l_returnflag_cmd_lastIdx,
      l_returnflag_cmd_tag         => PriceSummary_inst_l_returnflag_cmd_tag,
      l_linestatus_cmd_valid       => PriceSummary_inst_l_linestatus_cmd_valid,
      l_linestatus_cmd_ready       => PriceSummary_inst_l_linestatus_cmd_ready,
      l_linestatus_cmd_firstIdx    => PriceSummary_inst_l_linestatus_cmd_firstIdx,
      l_linestatus_cmd_lastIdx     => PriceSummary_inst_l_linestatus_cmd_lastIdx,
      l_linestatus_cmd_tag         => PriceSummary_inst_l_linestatus_cmd_tag,
      l_shipdate_cmd_valid         => PriceSummary_inst_l_shipdate_cmd_valid,
      l_shipdate_cmd_ready         => PriceSummary_inst_l_shipdate_cmd_ready,
      l_shipdate_cmd_firstIdx      => PriceSummary_inst_l_shipdate_cmd_firstIdx,
      l_shipdate_cmd_lastIdx       => PriceSummary_inst_l_shipdate_cmd_lastIdx,
      l_shipdate_cmd_tag           => PriceSummary_inst_l_shipdate_cmd_tag,
      start                        => PriceSummary_inst_start,
      stop                         => PriceSummary_inst_stop,
      reset                        => PriceSummary_inst_reset,
      idle                         => PriceSummary_inst_idle,
      busy                         => PriceSummary_inst_busy,
      done                         => PriceSummary_inst_done,
      result                       => PriceSummary_inst_result,
      l_firstidx                   => PriceSummary_inst_l_firstidx,
      l_lastidx                    => PriceSummary_inst_l_lastidx,
      rhigh                        => PriceSummary_inst_rhigh,
      rlow                         => PriceSummary_inst_rlow,
      status_1                     => PriceSummary_inst_status_1,
      status_2                     => PriceSummary_inst_status_2,
      r1                           => PriceSummary_inst_r1,
      r2                           => PriceSummary_inst_r2,
      r3                           => PriceSummary_inst_r3,
      r4                           => PriceSummary_inst_r4,
      r5                           => PriceSummary_inst_r5,
      r6                           => PriceSummary_inst_r6,
      r7                           => PriceSummary_inst_r7,
      r8                           => PriceSummary_inst_r8
    );

  mmio_inst : mmio
    port map (
      kcd_clk                       => kcd_clk,
      kcd_reset                     => kcd_reset,
      f_start_data                  => mmio_inst_f_start_data,
      f_stop_data                   => mmio_inst_f_stop_data,
      f_reset_data                  => mmio_inst_f_reset_data,
      f_idle_write_data             => mmio_inst_f_idle_write_data,
      f_busy_write_data             => mmio_inst_f_busy_write_data,
      f_done_write_data             => mmio_inst_f_done_write_data,
      f_result_write_data           => mmio_inst_f_result_write_data,
      f_l_firstidx_data             => mmio_inst_f_l_firstidx_data,
      f_l_lastidx_data              => mmio_inst_f_l_lastidx_data,
      f_l_quantity_values_data      => mmio_inst_f_l_quantity_values_data,
      f_l_extendedprice_values_data => mmio_inst_f_l_extendedprice_values_data,
      f_l_discount_values_data      => mmio_inst_f_l_discount_values_data,
      f_l_tax_values_data           => mmio_inst_f_l_tax_values_data,
      f_l_returnflag_offsets_data   => mmio_inst_f_l_returnflag_offsets_data,
      f_l_returnflag_values_data    => mmio_inst_f_l_returnflag_values_data,
      f_l_linestatus_offsets_data   => mmio_inst_f_l_linestatus_offsets_data,
      f_l_linestatus_values_data    => mmio_inst_f_l_linestatus_values_data,
      f_l_shipdate_values_data      => mmio_inst_f_l_shipdate_values_data,
      f_rhigh_write_data            => mmio_inst_f_rhigh_write_data,
      f_rlow_write_data             => mmio_inst_f_rlow_write_data,
      f_status_1_write_data         => mmio_inst_f_status_1_write_data,
      f_status_2_write_data         => mmio_inst_f_status_2_write_data,
      f_r1_write_data               => mmio_inst_f_r1_write_data,
      f_r2_write_data               => mmio_inst_f_r2_write_data,
      f_r3_write_data               => mmio_inst_f_r3_write_data,
      f_r4_write_data               => mmio_inst_f_r4_write_data,
      f_r5_write_data               => mmio_inst_f_r5_write_data,
      f_r6_write_data               => mmio_inst_f_r6_write_data,
      f_r7_write_data               => mmio_inst_f_r7_write_data,
      f_r8_write_data               => mmio_inst_f_r8_write_data,
      mmio_awvalid                  => mmio_inst_mmio_awvalid,
      mmio_awready                  => mmio_inst_mmio_awready,
      mmio_awaddr                   => mmio_inst_mmio_awaddr,
      mmio_wvalid                   => mmio_inst_mmio_wvalid,
      mmio_wready                   => mmio_inst_mmio_wready,
      mmio_wdata                    => mmio_inst_mmio_wdata,
      mmio_wstrb                    => mmio_inst_mmio_wstrb,
      mmio_bvalid                   => mmio_inst_mmio_bvalid,
      mmio_bready                   => mmio_inst_mmio_bready,
      mmio_bresp                    => mmio_inst_mmio_bresp,
      mmio_arvalid                  => mmio_inst_mmio_arvalid,
      mmio_arready                  => mmio_inst_mmio_arready,
      mmio_araddr                   => mmio_inst_mmio_araddr,
      mmio_rvalid                   => mmio_inst_mmio_rvalid,
      mmio_rready                   => mmio_inst_mmio_rready,
      mmio_rdata                    => mmio_inst_mmio_rdata,
      mmio_rresp                    => mmio_inst_mmio_rresp
    );

  l_quantity_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => L_QUANTITY_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => l_quantity_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => l_quantity_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => l_quantity_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => l_quantity_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => l_quantity_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => l_quantity_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => l_quantity_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => l_quantity_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => l_quantity_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => l_quantity_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => l_quantity_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => l_quantity_cmd_accm_inst_ctrl
    );

  l_extendedprice_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => L_EXTENDEDPRICE_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => l_extendedprice_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => l_extendedprice_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => l_extendedprice_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => l_extendedprice_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => l_extendedprice_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => l_extendedprice_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => l_extendedprice_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => l_extendedprice_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => l_extendedprice_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => l_extendedprice_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => l_extendedprice_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => l_extendedprice_cmd_accm_inst_ctrl
    );

  l_discount_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => L_DISCOUNT_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => l_discount_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => l_discount_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => l_discount_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => l_discount_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => l_discount_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => l_discount_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => l_discount_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => l_discount_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => l_discount_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => l_discount_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => l_discount_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => l_discount_cmd_accm_inst_ctrl
    );

  l_tax_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => L_TAX_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => l_tax_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => l_tax_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => l_tax_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => l_tax_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => l_tax_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => l_tax_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => l_tax_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => l_tax_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => l_tax_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => l_tax_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => l_tax_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => l_tax_cmd_accm_inst_ctrl
    );

  l_returnflag_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 2,
      BUS_ADDR_WIDTH => L_RETURNFLAG_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => l_returnflag_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => l_returnflag_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => l_returnflag_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => l_returnflag_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => l_returnflag_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => l_returnflag_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => l_returnflag_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => l_returnflag_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => l_returnflag_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => l_returnflag_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => l_returnflag_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => l_returnflag_cmd_accm_inst_ctrl
    );

  l_linestatus_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 2,
      BUS_ADDR_WIDTH => L_LINESTATUS_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => l_linestatus_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => l_linestatus_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => l_linestatus_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => l_linestatus_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => l_linestatus_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => l_linestatus_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => l_linestatus_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => l_linestatus_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => l_linestatus_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => l_linestatus_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => l_linestatus_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => l_linestatus_cmd_accm_inst_ctrl
    );

  l_shipdate_cmd_accm_inst : ArrayCmdCtrlMerger
    generic map (
      NUM_ADDR       => 1,
      BUS_ADDR_WIDTH => L_SHIPDATE_BUS_ADDR_WIDTH,
      INDEX_WIDTH    => INDEX_WIDTH,
      TAG_WIDTH      => TAG_WIDTH
    )
    port map (
      kernel_cmd_valid     => l_shipdate_cmd_accm_inst_kernel_cmd_valid,
      kernel_cmd_ready     => l_shipdate_cmd_accm_inst_kernel_cmd_ready,
      kernel_cmd_firstIdx  => l_shipdate_cmd_accm_inst_kernel_cmd_firstIdx,
      kernel_cmd_lastIdx   => l_shipdate_cmd_accm_inst_kernel_cmd_lastIdx,
      kernel_cmd_tag       => l_shipdate_cmd_accm_inst_kernel_cmd_tag,
      nucleus_cmd_valid    => l_shipdate_cmd_accm_inst_nucleus_cmd_valid,
      nucleus_cmd_ready    => l_shipdate_cmd_accm_inst_nucleus_cmd_ready,
      nucleus_cmd_firstIdx => l_shipdate_cmd_accm_inst_nucleus_cmd_firstIdx,
      nucleus_cmd_lastIdx  => l_shipdate_cmd_accm_inst_nucleus_cmd_lastIdx,
      nucleus_cmd_ctrl     => l_shipdate_cmd_accm_inst_nucleus_cmd_ctrl,
      nucleus_cmd_tag      => l_shipdate_cmd_accm_inst_nucleus_cmd_tag,
      ctrl                 => l_shipdate_cmd_accm_inst_ctrl
    );

  l_quantity_cmd_valid                            <= l_quantity_cmd_accm_inst_nucleus_cmd_valid;
  l_quantity_cmd_accm_inst_nucleus_cmd_ready      <= l_quantity_cmd_ready;
  l_quantity_cmd_firstIdx                         <= l_quantity_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_quantity_cmd_lastIdx                          <= l_quantity_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_quantity_cmd_ctrl                             <= l_quantity_cmd_accm_inst_nucleus_cmd_ctrl;
  l_quantity_cmd_tag                              <= l_quantity_cmd_accm_inst_nucleus_cmd_tag;

  l_extendedprice_cmd_valid                       <= l_extendedprice_cmd_accm_inst_nucleus_cmd_valid;
  l_extendedprice_cmd_accm_inst_nucleus_cmd_ready <= l_extendedprice_cmd_ready;
  l_extendedprice_cmd_firstIdx                    <= l_extendedprice_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_extendedprice_cmd_lastIdx                     <= l_extendedprice_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_extendedprice_cmd_ctrl                        <= l_extendedprice_cmd_accm_inst_nucleus_cmd_ctrl;
  l_extendedprice_cmd_tag                         <= l_extendedprice_cmd_accm_inst_nucleus_cmd_tag;

  l_discount_cmd_valid                            <= l_discount_cmd_accm_inst_nucleus_cmd_valid;
  l_discount_cmd_accm_inst_nucleus_cmd_ready      <= l_discount_cmd_ready;
  l_discount_cmd_firstIdx                         <= l_discount_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_discount_cmd_lastIdx                          <= l_discount_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_discount_cmd_ctrl                             <= l_discount_cmd_accm_inst_nucleus_cmd_ctrl;
  l_discount_cmd_tag                              <= l_discount_cmd_accm_inst_nucleus_cmd_tag;

  l_tax_cmd_valid                                 <= l_tax_cmd_accm_inst_nucleus_cmd_valid;
  l_tax_cmd_accm_inst_nucleus_cmd_ready           <= l_tax_cmd_ready;
  l_tax_cmd_firstIdx                              <= l_tax_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_tax_cmd_lastIdx                               <= l_tax_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_tax_cmd_ctrl                                  <= l_tax_cmd_accm_inst_nucleus_cmd_ctrl;
  l_tax_cmd_tag                                   <= l_tax_cmd_accm_inst_nucleus_cmd_tag;

  l_returnflag_cmd_valid                          <= l_returnflag_cmd_accm_inst_nucleus_cmd_valid;
  l_returnflag_cmd_accm_inst_nucleus_cmd_ready    <= l_returnflag_cmd_ready;
  l_returnflag_cmd_firstIdx                       <= l_returnflag_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_returnflag_cmd_lastIdx                        <= l_returnflag_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_returnflag_cmd_ctrl                           <= l_returnflag_cmd_accm_inst_nucleus_cmd_ctrl;
  l_returnflag_cmd_tag                            <= l_returnflag_cmd_accm_inst_nucleus_cmd_tag;

  l_linestatus_cmd_valid                          <= l_linestatus_cmd_accm_inst_nucleus_cmd_valid;
  l_linestatus_cmd_accm_inst_nucleus_cmd_ready    <= l_linestatus_cmd_ready;
  l_linestatus_cmd_firstIdx                       <= l_linestatus_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_linestatus_cmd_lastIdx                        <= l_linestatus_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_linestatus_cmd_ctrl                           <= l_linestatus_cmd_accm_inst_nucleus_cmd_ctrl;
  l_linestatus_cmd_tag                            <= l_linestatus_cmd_accm_inst_nucleus_cmd_tag;

  l_shipdate_cmd_valid                            <= l_shipdate_cmd_accm_inst_nucleus_cmd_valid;
  l_shipdate_cmd_accm_inst_nucleus_cmd_ready      <= l_shipdate_cmd_ready;
  l_shipdate_cmd_firstIdx                         <= l_shipdate_cmd_accm_inst_nucleus_cmd_firstIdx;
  l_shipdate_cmd_lastIdx                          <= l_shipdate_cmd_accm_inst_nucleus_cmd_lastIdx;
  l_shipdate_cmd_ctrl                             <= l_shipdate_cmd_accm_inst_nucleus_cmd_ctrl;
  l_shipdate_cmd_tag                              <= l_shipdate_cmd_accm_inst_nucleus_cmd_tag;

  PriceSummary_inst_l_quantity_valid                <= l_quantity_valid;
  l_quantity_ready                                  <= PriceSummary_inst_l_quantity_ready;
  PriceSummary_inst_l_quantity_dvalid               <= l_quantity_dvalid;
  PriceSummary_inst_l_quantity_last                 <= l_quantity_last;
  PriceSummary_inst_l_quantity                      <= l_quantity;

  PriceSummary_inst_l_extendedprice_valid           <= l_extendedprice_valid;
  l_extendedprice_ready                             <= PriceSummary_inst_l_extendedprice_ready;
  PriceSummary_inst_l_extendedprice_dvalid          <= l_extendedprice_dvalid;
  PriceSummary_inst_l_extendedprice_last            <= l_extendedprice_last;
  PriceSummary_inst_l_extendedprice                 <= l_extendedprice;

  PriceSummary_inst_l_discount_valid                <= l_discount_valid;
  l_discount_ready                                  <= PriceSummary_inst_l_discount_ready;
  PriceSummary_inst_l_discount_dvalid               <= l_discount_dvalid;
  PriceSummary_inst_l_discount_last                 <= l_discount_last;
  PriceSummary_inst_l_discount                      <= l_discount;

  PriceSummary_inst_l_tax_valid                     <= l_tax_valid;
  l_tax_ready                                       <= PriceSummary_inst_l_tax_ready;
  PriceSummary_inst_l_tax_dvalid                    <= l_tax_dvalid;
  PriceSummary_inst_l_tax_last                      <= l_tax_last;
  PriceSummary_inst_l_tax                           <= l_tax;

  PriceSummary_inst_l_returnflag_valid              <= l_returnflag_valid;
  l_returnflag_ready                                <= PriceSummary_inst_l_returnflag_ready;
  PriceSummary_inst_l_returnflag_dvalid             <= l_returnflag_dvalid;
  PriceSummary_inst_l_returnflag_last               <= l_returnflag_last;
  PriceSummary_inst_l_returnflag_length             <= l_returnflag_length;
  PriceSummary_inst_l_returnflag_count              <= l_returnflag_count;
  PriceSummary_inst_l_returnflag_chars_valid        <= l_returnflag_chars_valid;
  l_returnflag_chars_ready                          <= PriceSummary_inst_l_returnflag_chars_ready;
  PriceSummary_inst_l_returnflag_chars_dvalid       <= l_returnflag_chars_dvalid;
  PriceSummary_inst_l_returnflag_chars_last         <= l_returnflag_chars_last;
  PriceSummary_inst_l_returnflag_chars              <= l_returnflag_chars;
  PriceSummary_inst_l_returnflag_chars_count        <= l_returnflag_chars_count;

  PriceSummary_inst_l_linestatus_valid              <= l_linestatus_valid;
  l_linestatus_ready                                <= PriceSummary_inst_l_linestatus_ready;
  PriceSummary_inst_l_linestatus_dvalid             <= l_linestatus_dvalid;
  PriceSummary_inst_l_linestatus_last               <= l_linestatus_last;
  PriceSummary_inst_l_linestatus_length             <= l_linestatus_length;
  PriceSummary_inst_l_linestatus_count              <= l_linestatus_count;
  PriceSummary_inst_l_linestatus_chars_valid        <= l_linestatus_chars_valid;
  l_linestatus_chars_ready                          <= PriceSummary_inst_l_linestatus_chars_ready;
  PriceSummary_inst_l_linestatus_chars_dvalid       <= l_linestatus_chars_dvalid;
  PriceSummary_inst_l_linestatus_chars_last         <= l_linestatus_chars_last;
  PriceSummary_inst_l_linestatus_chars              <= l_linestatus_chars;
  PriceSummary_inst_l_linestatus_chars_count        <= l_linestatus_chars_count;

  PriceSummary_inst_l_shipdate_valid                <= l_shipdate_valid;
  l_shipdate_ready                                  <= PriceSummary_inst_l_shipdate_ready;
  PriceSummary_inst_l_shipdate_dvalid               <= l_shipdate_dvalid;
  PriceSummary_inst_l_shipdate_last                 <= l_shipdate_last;
  PriceSummary_inst_l_shipdate                      <= l_shipdate;

  PriceSummary_inst_l_quantity_unl_valid            <= l_quantity_unl_valid;
  l_quantity_unl_ready                              <= PriceSummary_inst_l_quantity_unl_ready;
  PriceSummary_inst_l_quantity_unl_tag              <= l_quantity_unl_tag;

  PriceSummary_inst_l_extendedprice_unl_valid       <= l_extendedprice_unl_valid;
  l_extendedprice_unl_ready                         <= PriceSummary_inst_l_extendedprice_unl_ready;
  PriceSummary_inst_l_extendedprice_unl_tag         <= l_extendedprice_unl_tag;

  PriceSummary_inst_l_discount_unl_valid            <= l_discount_unl_valid;
  l_discount_unl_ready                              <= PriceSummary_inst_l_discount_unl_ready;
  PriceSummary_inst_l_discount_unl_tag              <= l_discount_unl_tag;

  PriceSummary_inst_l_tax_unl_valid                 <= l_tax_unl_valid;
  l_tax_unl_ready                                   <= PriceSummary_inst_l_tax_unl_ready;
  PriceSummary_inst_l_tax_unl_tag                   <= l_tax_unl_tag;

  PriceSummary_inst_l_returnflag_unl_valid          <= l_returnflag_unl_valid;
  l_returnflag_unl_ready                            <= PriceSummary_inst_l_returnflag_unl_ready;
  PriceSummary_inst_l_returnflag_unl_tag            <= l_returnflag_unl_tag;

  PriceSummary_inst_l_linestatus_unl_valid          <= l_linestatus_unl_valid;
  l_linestatus_unl_ready                            <= PriceSummary_inst_l_linestatus_unl_ready;
  PriceSummary_inst_l_linestatus_unl_tag            <= l_linestatus_unl_tag;

  PriceSummary_inst_l_shipdate_unl_valid            <= l_shipdate_unl_valid;
  l_shipdate_unl_ready                              <= PriceSummary_inst_l_shipdate_unl_ready;
  PriceSummary_inst_l_shipdate_unl_tag              <= l_shipdate_unl_tag;

  PriceSummary_inst_start                           <= mmio_inst_f_start_data;
  PriceSummary_inst_stop                            <= mmio_inst_f_stop_data;
  PriceSummary_inst_reset                           <= mmio_inst_f_reset_data;
  PriceSummary_inst_l_firstidx                      <= mmio_inst_f_l_firstidx_data;
  PriceSummary_inst_l_lastidx                       <= mmio_inst_f_l_lastidx_data;
  mmio_inst_f_idle_write_data                       <= PriceSummary_inst_idle;
  mmio_inst_f_busy_write_data                       <= PriceSummary_inst_busy;
  mmio_inst_f_done_write_data                       <= PriceSummary_inst_done;
  mmio_inst_f_result_write_data                     <= PriceSummary_inst_result;
  mmio_inst_f_rhigh_write_data                      <= PriceSummary_inst_rhigh;
  mmio_inst_f_rlow_write_data                       <= PriceSummary_inst_rlow;
  mmio_inst_f_status_1_write_data                   <= PriceSummary_inst_status_1;
  mmio_inst_f_status_2_write_data                   <= PriceSummary_inst_status_2;
  mmio_inst_f_r1_write_data                         <= PriceSummary_inst_r1;
  mmio_inst_f_r2_write_data                         <= PriceSummary_inst_r2;
  mmio_inst_f_r3_write_data                         <= PriceSummary_inst_r3;
  mmio_inst_f_r4_write_data                         <= PriceSummary_inst_r4;
  mmio_inst_f_r5_write_data                         <= PriceSummary_inst_r5;
  mmio_inst_f_r6_write_data                         <= PriceSummary_inst_r6;
  mmio_inst_f_r7_write_data                         <= PriceSummary_inst_r7;
  mmio_inst_f_r8_write_data                         <= PriceSummary_inst_r8;
  mmio_inst_mmio_awvalid                            <= mmio_awvalid;
  mmio_awready                                      <= mmio_inst_mmio_awready;
  mmio_inst_mmio_awaddr                             <= mmio_awaddr;
  mmio_inst_mmio_wvalid                             <= mmio_wvalid;
  mmio_wready                                       <= mmio_inst_mmio_wready;
  mmio_inst_mmio_wdata                              <= mmio_wdata;
  mmio_inst_mmio_wstrb                              <= mmio_wstrb;
  mmio_bvalid                                       <= mmio_inst_mmio_bvalid;
  mmio_inst_mmio_bready                             <= mmio_bready;
  mmio_bresp                                        <= mmio_inst_mmio_bresp;
  mmio_inst_mmio_arvalid                            <= mmio_arvalid;
  mmio_arready                                      <= mmio_inst_mmio_arready;
  mmio_inst_mmio_araddr                             <= mmio_araddr;
  mmio_rvalid                                       <= mmio_inst_mmio_rvalid;
  mmio_inst_mmio_rready                             <= mmio_rready;
  mmio_rdata                                        <= mmio_inst_mmio_rdata;
  mmio_rresp                                        <= mmio_inst_mmio_rresp;

  l_quantity_cmd_accm_inst_kernel_cmd_valid         <= PriceSummary_inst_l_quantity_cmd_valid;
  PriceSummary_inst_l_quantity_cmd_ready            <= l_quantity_cmd_accm_inst_kernel_cmd_ready;
  l_quantity_cmd_accm_inst_kernel_cmd_firstIdx      <= PriceSummary_inst_l_quantity_cmd_firstIdx;
  l_quantity_cmd_accm_inst_kernel_cmd_lastIdx       <= PriceSummary_inst_l_quantity_cmd_lastIdx;
  l_quantity_cmd_accm_inst_kernel_cmd_tag           <= PriceSummary_inst_l_quantity_cmd_tag;

  l_extendedprice_cmd_accm_inst_kernel_cmd_valid    <= PriceSummary_inst_l_extendedprice_cmd_valid;
  PriceSummary_inst_l_extendedprice_cmd_ready       <= l_extendedprice_cmd_accm_inst_kernel_cmd_ready;
  l_extendedprice_cmd_accm_inst_kernel_cmd_firstIdx <= PriceSummary_inst_l_extendedprice_cmd_firstIdx;
  l_extendedprice_cmd_accm_inst_kernel_cmd_lastIdx  <= PriceSummary_inst_l_extendedprice_cmd_lastIdx;
  l_extendedprice_cmd_accm_inst_kernel_cmd_tag      <= PriceSummary_inst_l_extendedprice_cmd_tag;

  l_discount_cmd_accm_inst_kernel_cmd_valid         <= PriceSummary_inst_l_discount_cmd_valid;
  PriceSummary_inst_l_discount_cmd_ready            <= l_discount_cmd_accm_inst_kernel_cmd_ready;
  l_discount_cmd_accm_inst_kernel_cmd_firstIdx      <= PriceSummary_inst_l_discount_cmd_firstIdx;
  l_discount_cmd_accm_inst_kernel_cmd_lastIdx       <= PriceSummary_inst_l_discount_cmd_lastIdx;
  l_discount_cmd_accm_inst_kernel_cmd_tag           <= PriceSummary_inst_l_discount_cmd_tag;

  l_tax_cmd_accm_inst_kernel_cmd_valid              <= PriceSummary_inst_l_tax_cmd_valid;
  PriceSummary_inst_l_tax_cmd_ready                 <= l_tax_cmd_accm_inst_kernel_cmd_ready;
  l_tax_cmd_accm_inst_kernel_cmd_firstIdx           <= PriceSummary_inst_l_tax_cmd_firstIdx;
  l_tax_cmd_accm_inst_kernel_cmd_lastIdx            <= PriceSummary_inst_l_tax_cmd_lastIdx;
  l_tax_cmd_accm_inst_kernel_cmd_tag                <= PriceSummary_inst_l_tax_cmd_tag;

  l_returnflag_cmd_accm_inst_kernel_cmd_valid       <= PriceSummary_inst_l_returnflag_cmd_valid;
  PriceSummary_inst_l_returnflag_cmd_ready          <= l_returnflag_cmd_accm_inst_kernel_cmd_ready;
  l_returnflag_cmd_accm_inst_kernel_cmd_firstIdx    <= PriceSummary_inst_l_returnflag_cmd_firstIdx;
  l_returnflag_cmd_accm_inst_kernel_cmd_lastIdx     <= PriceSummary_inst_l_returnflag_cmd_lastIdx;
  l_returnflag_cmd_accm_inst_kernel_cmd_tag         <= PriceSummary_inst_l_returnflag_cmd_tag;

  l_linestatus_cmd_accm_inst_kernel_cmd_valid       <= PriceSummary_inst_l_linestatus_cmd_valid;
  PriceSummary_inst_l_linestatus_cmd_ready          <= l_linestatus_cmd_accm_inst_kernel_cmd_ready;
  l_linestatus_cmd_accm_inst_kernel_cmd_firstIdx    <= PriceSummary_inst_l_linestatus_cmd_firstIdx;
  l_linestatus_cmd_accm_inst_kernel_cmd_lastIdx     <= PriceSummary_inst_l_linestatus_cmd_lastIdx;
  l_linestatus_cmd_accm_inst_kernel_cmd_tag         <= PriceSummary_inst_l_linestatus_cmd_tag;

  l_shipdate_cmd_accm_inst_kernel_cmd_valid         <= PriceSummary_inst_l_shipdate_cmd_valid;
  PriceSummary_inst_l_shipdate_cmd_ready            <= l_shipdate_cmd_accm_inst_kernel_cmd_ready;
  l_shipdate_cmd_accm_inst_kernel_cmd_firstIdx      <= PriceSummary_inst_l_shipdate_cmd_firstIdx;
  l_shipdate_cmd_accm_inst_kernel_cmd_lastIdx       <= PriceSummary_inst_l_shipdate_cmd_lastIdx;
  l_shipdate_cmd_accm_inst_kernel_cmd_tag           <= PriceSummary_inst_l_shipdate_cmd_tag;

  l_quantity_cmd_accm_inst_ctrl(63 downto 0)      <= mmio_inst_f_l_quantity_values_data;
  l_extendedprice_cmd_accm_inst_ctrl(63 downto 0) <= mmio_inst_f_l_extendedprice_values_data;
  l_discount_cmd_accm_inst_ctrl(63 downto 0)      <= mmio_inst_f_l_discount_values_data;
  l_tax_cmd_accm_inst_ctrl(63 downto 0)           <= mmio_inst_f_l_tax_values_data;
  l_returnflag_cmd_accm_inst_ctrl(63 downto 0)    <= mmio_inst_f_l_returnflag_offsets_data;
  l_returnflag_cmd_accm_inst_ctrl(127 downto 64)  <= mmio_inst_f_l_returnflag_values_data;

  l_linestatus_cmd_accm_inst_ctrl(63 downto 0)    <= mmio_inst_f_l_linestatus_offsets_data;
  l_linestatus_cmd_accm_inst_ctrl(127 downto 64)  <= mmio_inst_f_l_linestatus_values_data;

  l_shipdate_cmd_accm_inst_ctrl(63 downto 0)      <= mmio_inst_f_l_shipdate_values_data;

end architecture;
