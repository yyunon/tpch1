-- Copyright 2018-2019 Delft University of Technology
--
-- Licensed under the Apache License, Version 2.0 (the "License");
-- you may not use this file except in compliance with the License.
-- You may obtain a copy of the License at
--
--     http://www.apache.org/licenses/LICENSE-2.0
--
-- Unless required by applicable law or agreed to in writing, software
-- distributed under the License is distributed on an "AS IS" BASIS,
-- WITHOUT WARRANTIES OR CONDITIONS OF ANY KIND, either express or implied.
-- See the License for the specific language governing permissions and
-- limitations under the License.
--
-- This file was generated by Fletchgen. Modify this file at your own risk.

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity PriceSummary is
  generic (
    INDEX_WIDTH : integer := 32;
    TAG_WIDTH   : integer := 1
  );
  port (
    kcd_clk                      : in  std_logic;
    kcd_reset                    : in  std_logic;
    l_quantity_valid             : in  std_logic;
    l_quantity_ready             : out std_logic;
    l_quantity_dvalid            : in  std_logic;
    l_quantity_last              : in  std_logic;
    l_quantity                   : in  std_logic_vector(63 downto 0);
    l_extendedprice_valid        : in  std_logic;
    l_extendedprice_ready        : out std_logic;
    l_extendedprice_dvalid       : in  std_logic;
    l_extendedprice_last         : in  std_logic;
    l_extendedprice              : in  std_logic_vector(63 downto 0);
    l_discount_valid             : in  std_logic;
    l_discount_ready             : out std_logic;
    l_discount_dvalid            : in  std_logic;
    l_discount_last              : in  std_logic;
    l_discount                   : in  std_logic_vector(63 downto 0);
    l_tax_valid                  : in  std_logic;
    l_tax_ready                  : out std_logic;
    l_tax_dvalid                 : in  std_logic;
    l_tax_last                   : in  std_logic;
    l_tax                        : in  std_logic_vector(63 downto 0);
    l_returnflag_valid           : in  std_logic;
    l_returnflag_ready           : out std_logic;
    l_returnflag_dvalid          : in  std_logic;
    l_returnflag_last            : in  std_logic;
    l_returnflag_length          : in  std_logic_vector(31 downto 0);
    l_returnflag_count           : in  std_logic_vector(0 downto 0);
    l_returnflag_chars_valid     : in  std_logic;
    l_returnflag_chars_ready     : out std_logic;
    l_returnflag_chars_dvalid    : in  std_logic;
    l_returnflag_chars_last      : in  std_logic;
    l_returnflag_chars           : in  std_logic_vector(7 downto 0);
    l_returnflag_chars_count     : in  std_logic_vector(0 downto 0);
    l_linestatus_valid           : in  std_logic;
    l_linestatus_ready           : out std_logic;
    l_linestatus_dvalid          : in  std_logic;
    l_linestatus_last            : in  std_logic;
    l_linestatus_length          : in  std_logic_vector(31 downto 0);
    l_linestatus_count           : in  std_logic_vector(0 downto 0);
    l_linestatus_chars_valid     : in  std_logic;
    l_linestatus_chars_ready     : out std_logic;
    l_linestatus_chars_dvalid    : in  std_logic;
    l_linestatus_chars_last      : in  std_logic;
    l_linestatus_chars           : in  std_logic_vector(7 downto 0);
    l_linestatus_chars_count     : in  std_logic_vector(0 downto 0);
    l_shipdate_valid             : in  std_logic;
    l_shipdate_ready             : out std_logic;
    l_shipdate_dvalid            : in  std_logic;
    l_shipdate_last              : in  std_logic;
    l_shipdate                   : in  std_logic_vector(31 downto 0);
    l_quantity_unl_valid         : in  std_logic;
    l_quantity_unl_ready         : out std_logic;
    l_quantity_unl_tag           : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_extendedprice_unl_valid    : in  std_logic;
    l_extendedprice_unl_ready    : out std_logic;
    l_extendedprice_unl_tag      : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_discount_unl_valid         : in  std_logic;
    l_discount_unl_ready         : out std_logic;
    l_discount_unl_tag           : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_tax_unl_valid              : in  std_logic;
    l_tax_unl_ready              : out std_logic;
    l_tax_unl_tag                : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_returnflag_unl_valid       : in  std_logic;
    l_returnflag_unl_ready       : out std_logic;
    l_returnflag_unl_tag         : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_linestatus_unl_valid       : in  std_logic;
    l_linestatus_unl_ready       : out std_logic;
    l_linestatus_unl_tag         : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_shipdate_unl_valid         : in  std_logic;
    l_shipdate_unl_ready         : out std_logic;
    l_shipdate_unl_tag           : in  std_logic_vector(TAG_WIDTH-1 downto 0);
    l_quantity_cmd_valid         : out std_logic;
    l_quantity_cmd_ready         : in  std_logic;
    l_quantity_cmd_firstIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_quantity_cmd_lastIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_quantity_cmd_tag           : out std_logic_vector(TAG_WIDTH-1 downto 0);
    l_extendedprice_cmd_valid    : out std_logic;
    l_extendedprice_cmd_ready    : in  std_logic;
    l_extendedprice_cmd_firstIdx : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_extendedprice_cmd_lastIdx  : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_extendedprice_cmd_tag      : out std_logic_vector(TAG_WIDTH-1 downto 0);
    l_discount_cmd_valid         : out std_logic;
    l_discount_cmd_ready         : in  std_logic;
    l_discount_cmd_firstIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_discount_cmd_lastIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_discount_cmd_tag           : out std_logic_vector(TAG_WIDTH-1 downto 0);
    l_tax_cmd_valid              : out std_logic;
    l_tax_cmd_ready              : in  std_logic;
    l_tax_cmd_firstIdx           : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_tax_cmd_lastIdx            : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_tax_cmd_tag                : out std_logic_vector(TAG_WIDTH-1 downto 0);
    l_returnflag_cmd_valid       : out std_logic;
    l_returnflag_cmd_ready       : in  std_logic;
    l_returnflag_cmd_firstIdx    : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_returnflag_cmd_lastIdx     : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_returnflag_cmd_tag         : out std_logic_vector(TAG_WIDTH-1 downto 0);
    l_linestatus_cmd_valid       : out std_logic;
    l_linestatus_cmd_ready       : in  std_logic;
    l_linestatus_cmd_firstIdx    : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_linestatus_cmd_lastIdx     : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_linestatus_cmd_tag         : out std_logic_vector(TAG_WIDTH-1 downto 0);
    l_shipdate_cmd_valid         : out std_logic;
    l_shipdate_cmd_ready         : in  std_logic;
    l_shipdate_cmd_firstIdx      : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_shipdate_cmd_lastIdx       : out std_logic_vector(INDEX_WIDTH-1 downto 0);
    l_shipdate_cmd_tag           : out std_logic_vector(TAG_WIDTH-1 downto 0);
    start                        : in  std_logic;
    stop                         : in  std_logic;
    reset                        : in  std_logic;
    idle                         : out std_logic;
    busy                         : out std_logic;
    done                         : out std_logic;
    result                       : out std_logic_vector(63 downto 0);
    l_firstidx                   : in  std_logic_vector(31 downto 0);
    l_lastidx                    : in  std_logic_vector(31 downto 0);
    rhigh                        : out std_logic_vector(31 downto 0);
    rlow                         : out std_logic_vector(31 downto 0);
    status_1                     : out std_logic_vector(31 downto 0);
    status_2                     : out std_logic_vector(31 downto 0);
    r1                           : out std_logic_vector(63 downto 0);
    r2                           : out std_logic_vector(63 downto 0);
    r3                           : out std_logic_vector(63 downto 0);
    r4                           : out std_logic_vector(63 downto 0);
    r5                           : out std_logic_vector(63 downto 0);
    r6                           : out std_logic_vector(63 downto 0);
    r7                           : out std_logic_vector(63 downto 0);
    r8                           : out std_logic_vector(63 downto 0)
  );
end entity;

architecture Implementation of PriceSummary is
begin
end architecture;
